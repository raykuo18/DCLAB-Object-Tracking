// w_r_idx
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };

// w_r_idx
