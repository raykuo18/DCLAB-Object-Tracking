// w_pos_ptr
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000011,
        `W_POS_PTR_BITWIDTH'b00000000110,
        `W_POS_PTR_BITWIDTH'b00000001001,
        `W_POS_PTR_BITWIDTH'b00000001100,
        `W_POS_PTR_BITWIDTH'b00000001111,
        `W_POS_PTR_BITWIDTH'b00000010010,
        `W_POS_PTR_BITWIDTH'b00000010101,
        `W_POS_PTR_BITWIDTH'b00000011000,
        `W_POS_PTR_BITWIDTH'b00000011011,
        `W_POS_PTR_BITWIDTH'b00000011110,
        `W_POS_PTR_BITWIDTH'b00000100001,
        `W_POS_PTR_BITWIDTH'b00000100100,
        `W_POS_PTR_BITWIDTH'b00000100110,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000101010,
        `W_POS_PTR_BITWIDTH'b00000101101,
        `W_POS_PTR_BITWIDTH'b00000110000,
        `W_POS_PTR_BITWIDTH'b00000110011,
        `W_POS_PTR_BITWIDTH'b00000110110,
        `W_POS_PTR_BITWIDTH'b00000111001,
        `W_POS_PTR_BITWIDTH'b00000111011,
        `W_POS_PTR_BITWIDTH'b00000111110,
        `W_POS_PTR_BITWIDTH'b00000111110
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00001000100,
        `W_POS_PTR_BITWIDTH'b00001000111,
        `W_POS_PTR_BITWIDTH'b00001001001,
        `W_POS_PTR_BITWIDTH'b00001001100,
        `W_POS_PTR_BITWIDTH'b00001001111,
        `W_POS_PTR_BITWIDTH'b00001010001,
        `W_POS_PTR_BITWIDTH'b00001010100,
        `W_POS_PTR_BITWIDTH'b00001010111,
        `W_POS_PTR_BITWIDTH'b00001011000,
        `W_POS_PTR_BITWIDTH'b00001011011,
        `W_POS_PTR_BITWIDTH'b00001011110,
        `W_POS_PTR_BITWIDTH'b00001100001,
        `W_POS_PTR_BITWIDTH'b00001100100,
        `W_POS_PTR_BITWIDTH'b00001100111,
        `W_POS_PTR_BITWIDTH'b00001101010,
        `W_POS_PTR_BITWIDTH'b00001101101,
        `W_POS_PTR_BITWIDTH'b00001110000,
        `W_POS_PTR_BITWIDTH'b00001110011,
        `W_POS_PTR_BITWIDTH'b00001110110,
        `W_POS_PTR_BITWIDTH'b00001111001,
        `W_POS_PTR_BITWIDTH'b00001111100,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010000010,
        `W_POS_PTR_BITWIDTH'b00010000010
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00010000110,
        `W_POS_PTR_BITWIDTH'b00010001001,
        `W_POS_PTR_BITWIDTH'b00010001010,
        `W_POS_PTR_BITWIDTH'b00010001100,
        `W_POS_PTR_BITWIDTH'b00010001111,
        `W_POS_PTR_BITWIDTH'b00010010001,
        `W_POS_PTR_BITWIDTH'b00010010100,
        `W_POS_PTR_BITWIDTH'b00010010111,
        `W_POS_PTR_BITWIDTH'b00010011010,
        `W_POS_PTR_BITWIDTH'b00010011100,
        `W_POS_PTR_BITWIDTH'b00010011111,
        `W_POS_PTR_BITWIDTH'b00010100010,
        `W_POS_PTR_BITWIDTH'b00010100101,
        `W_POS_PTR_BITWIDTH'b00010100110,
        `W_POS_PTR_BITWIDTH'b00010101000,
        `W_POS_PTR_BITWIDTH'b00010101001,
        `W_POS_PTR_BITWIDTH'b00010101100,
        `W_POS_PTR_BITWIDTH'b00010101111,
        `W_POS_PTR_BITWIDTH'b00010110010,
        `W_POS_PTR_BITWIDTH'b00010110101,
        `W_POS_PTR_BITWIDTH'b00010110110,
        `W_POS_PTR_BITWIDTH'b00010111001,
        `W_POS_PTR_BITWIDTH'b00010111100,
        `W_POS_PTR_BITWIDTH'b00010111100
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000010,
        `W_POS_PTR_BITWIDTH'b00000000110,
        `W_POS_PTR_BITWIDTH'b00000001010,
        `W_POS_PTR_BITWIDTH'b00000001100,
        `W_POS_PTR_BITWIDTH'b00000010000,
        `W_POS_PTR_BITWIDTH'b00000010011,
        `W_POS_PTR_BITWIDTH'b00000010100,
        `W_POS_PTR_BITWIDTH'b00000011001,
        `W_POS_PTR_BITWIDTH'b00000011100,
        `W_POS_PTR_BITWIDTH'b00000011111,
        `W_POS_PTR_BITWIDTH'b00000100010,
        `W_POS_PTR_BITWIDTH'b00000100101,
        `W_POS_PTR_BITWIDTH'b00000100111,
        `W_POS_PTR_BITWIDTH'b00000101100,
        `W_POS_PTR_BITWIDTH'b00000110001,
        `W_POS_PTR_BITWIDTH'b00000110101,
        `W_POS_PTR_BITWIDTH'b00000110111,
        `W_POS_PTR_BITWIDTH'b00000111001,
        `W_POS_PTR_BITWIDTH'b00000111110,
        `W_POS_PTR_BITWIDTH'b00001000001,
        `W_POS_PTR_BITWIDTH'b00001000100,
        `W_POS_PTR_BITWIDTH'b00001000110,
        `W_POS_PTR_BITWIDTH'b00001000110
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00001001110,
        `W_POS_PTR_BITWIDTH'b00001010011,
        `W_POS_PTR_BITWIDTH'b00001011000,
        `W_POS_PTR_BITWIDTH'b00001011010,
        `W_POS_PTR_BITWIDTH'b00001011101,
        `W_POS_PTR_BITWIDTH'b00001011111,
        `W_POS_PTR_BITWIDTH'b00001100010,
        `W_POS_PTR_BITWIDTH'b00001100110,
        `W_POS_PTR_BITWIDTH'b00001101010,
        `W_POS_PTR_BITWIDTH'b00001101110,
        `W_POS_PTR_BITWIDTH'b00001110001,
        `W_POS_PTR_BITWIDTH'b00001110100,
        `W_POS_PTR_BITWIDTH'b00001111001,
        `W_POS_PTR_BITWIDTH'b00001111101,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010000010,
        `W_POS_PTR_BITWIDTH'b00010000011,
        `W_POS_PTR_BITWIDTH'b00010001001,
        `W_POS_PTR_BITWIDTH'b00010001110,
        `W_POS_PTR_BITWIDTH'b00010010010,
        `W_POS_PTR_BITWIDTH'b00010010111,
        `W_POS_PTR_BITWIDTH'b00010011100,
        `W_POS_PTR_BITWIDTH'b00010011100
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00010100100,
        `W_POS_PTR_BITWIDTH'b00010101001,
        `W_POS_PTR_BITWIDTH'b00010101110,
        `W_POS_PTR_BITWIDTH'b00010110001,
        `W_POS_PTR_BITWIDTH'b00010110011,
        `W_POS_PTR_BITWIDTH'b00010111000,
        `W_POS_PTR_BITWIDTH'b00010111010,
        `W_POS_PTR_BITWIDTH'b00010111101,
        `W_POS_PTR_BITWIDTH'b00011000000,
        `W_POS_PTR_BITWIDTH'b00011000010,
        `W_POS_PTR_BITWIDTH'b00011000011,
        `W_POS_PTR_BITWIDTH'b00011001000,
        `W_POS_PTR_BITWIDTH'b00011001010,
        `W_POS_PTR_BITWIDTH'b00011001111,
        `W_POS_PTR_BITWIDTH'b00011010001,
        `W_POS_PTR_BITWIDTH'b00011010011,
        `W_POS_PTR_BITWIDTH'b00011010110,
        `W_POS_PTR_BITWIDTH'b00011010111,
        `W_POS_PTR_BITWIDTH'b00011011010,
        `W_POS_PTR_BITWIDTH'b00011011101,
        `W_POS_PTR_BITWIDTH'b00011100001,
        `W_POS_PTR_BITWIDTH'b00011100010,
        `W_POS_PTR_BITWIDTH'b00011100010
    };

// w_pos_ptr
