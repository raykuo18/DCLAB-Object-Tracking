// w_data
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_DATA_BITWIDTH'b1111110011100101,
        `W_DATA_BITWIDTH'b1111111001011110,
        `W_DATA_BITWIDTH'b0000001001011101,
        `W_DATA_BITWIDTH'b1111111101011000,
        `W_DATA_BITWIDTH'b1111110101101101,
        `W_DATA_BITWIDTH'b1111110010110110,
        `W_DATA_BITWIDTH'b0000001110111010,
        `W_DATA_BITWIDTH'b1111111010001100,
        `W_DATA_BITWIDTH'b0000001000001011,
        `W_DATA_BITWIDTH'b1111101111110111,
        `W_DATA_BITWIDTH'b0000000010111010,
        `W_DATA_BITWIDTH'b0000001101011100,
        `W_DATA_BITWIDTH'b0000000110001011,
        `W_DATA_BITWIDTH'b1111110000101100,
        `W_DATA_BITWIDTH'b0000001110000100,
        `W_DATA_BITWIDTH'b0000010011010001,
        `W_DATA_BITWIDTH'b1111100001100110,
        `W_DATA_BITWIDTH'b0000001110000111,
        `W_DATA_BITWIDTH'b1111110110101001,
        `W_DATA_BITWIDTH'b1111111000011000,
        `W_DATA_BITWIDTH'b0000001000010001,
        `W_DATA_BITWIDTH'b0000000110110111,
        `W_DATA_BITWIDTH'b0000000010000000,
        `W_DATA_BITWIDTH'b1111110100000000,
        `W_DATA_BITWIDTH'b0000000110010101,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b0000000101011011,
        `W_DATA_BITWIDTH'b0000001000101100,
        `W_DATA_BITWIDTH'b0000000111010100,
        `W_DATA_BITWIDTH'b1111111000001000,
        `W_DATA_BITWIDTH'b1111111011011010,
        `W_DATA_BITWIDTH'b0000000010011110,
        `W_DATA_BITWIDTH'b1111111100110001,
        `W_DATA_BITWIDTH'b0000010000101111,
        `W_DATA_BITWIDTH'b1111101001000011,
        `W_DATA_BITWIDTH'b1111111000011101,
        `W_DATA_BITWIDTH'b1111110010111111,
        `W_DATA_BITWIDTH'b1111111101110010,
        `W_DATA_BITWIDTH'b1111111011110001,
        `W_DATA_BITWIDTH'b1111111011100011,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000111100110,
        `W_DATA_BITWIDTH'b0000010001100000,
        `W_DATA_BITWIDTH'b1111101101100010,
        `W_DATA_BITWIDTH'b1111111101110110,
        `W_DATA_BITWIDTH'b0000001110000101,
        `W_DATA_BITWIDTH'b1111100111001110,
        `W_DATA_BITWIDTH'b0000000101011000,
        `W_DATA_BITWIDTH'b0000001101011101,
        `W_DATA_BITWIDTH'b1111110000000010,
        `W_DATA_BITWIDTH'b0000001000001000,
        `W_DATA_BITWIDTH'b1111100111110100,
        `W_DATA_BITWIDTH'b0000000111100011,
        `W_DATA_BITWIDTH'b0000001001010101,
        `W_DATA_BITWIDTH'b0000000100011010,
        `W_DATA_BITWIDTH'b0000010011000111,
        `W_DATA_BITWIDTH'b0000000010000001,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000000011100001,
        `W_DATA_BITWIDTH'b1111111010100101,
        `W_DATA_BITWIDTH'b0000000101001001,
        `W_DATA_BITWIDTH'b0000001111100110,
        `W_DATA_BITWIDTH'b0000001010101001,
        `W_DATA_BITWIDTH'b0000011011010011,
        `W_DATA_BITWIDTH'b1111101100010100,
        `W_DATA_BITWIDTH'b0000000010010101,
        `W_DATA_BITWIDTH'b1111101001100110,
        `W_DATA_BITWIDTH'b1111101001100110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_DATA_BITWIDTH'b0000001011111110,
        `W_DATA_BITWIDTH'b0000000001111100,
        `W_DATA_BITWIDTH'b0000000100001101,
        `W_DATA_BITWIDTH'b0000001001111011,
        `W_DATA_BITWIDTH'b1111111011100110,
        `W_DATA_BITWIDTH'b1111111010000111,
        `W_DATA_BITWIDTH'b1111101111000001,
        `W_DATA_BITWIDTH'b1111111101100001,
        `W_DATA_BITWIDTH'b0000011011100110,
        `W_DATA_BITWIDTH'b0000000011100101,
        `W_DATA_BITWIDTH'b1111110011101111,
        `W_DATA_BITWIDTH'b0000000011101000,
        `W_DATA_BITWIDTH'b1111110100010101,
        `W_DATA_BITWIDTH'b1111110010010100,
        `W_DATA_BITWIDTH'b1111110011100001,
        `W_DATA_BITWIDTH'b0000000101010100,
        `W_DATA_BITWIDTH'b1111110111011100,
        `W_DATA_BITWIDTH'b1111110111011000,
        `W_DATA_BITWIDTH'b0000000101001100,
        `W_DATA_BITWIDTH'b1111110100010011,
        `W_DATA_BITWIDTH'b1111111010011111,
        `W_DATA_BITWIDTH'b0000001001100101,
        `W_DATA_BITWIDTH'b0000000111010101,
        `W_DATA_BITWIDTH'b1111100101110011,
        `W_DATA_BITWIDTH'b0000011010010111,
        `W_DATA_BITWIDTH'b0000000011000011,
        `W_DATA_BITWIDTH'b1111110101101010,
        `W_DATA_BITWIDTH'b0000000110111011,
        `W_DATA_BITWIDTH'b1111101110111011,
        `W_DATA_BITWIDTH'b0000010111100100,
        `W_DATA_BITWIDTH'b0000000110001111,
        `W_DATA_BITWIDTH'b0000010000001011,
        `W_DATA_BITWIDTH'b1111110111001100,
        `W_DATA_BITWIDTH'b1111111001100010,
        `W_DATA_BITWIDTH'b0000000101110101,
        `W_DATA_BITWIDTH'b1111101101101110,
        `W_DATA_BITWIDTH'b0000000100001110,
        `W_DATA_BITWIDTH'b0000000110111001,
        `W_DATA_BITWIDTH'b1111111100110110,
        `W_DATA_BITWIDTH'b1111111100101010,
        `W_DATA_BITWIDTH'b0000000111111111,
        `W_DATA_BITWIDTH'b0000100101101101,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110000000101,
        `W_DATA_BITWIDTH'b1111110000011011,
        `W_DATA_BITWIDTH'b0000000010110101,
        `W_DATA_BITWIDTH'b0000011010110011,
        `W_DATA_BITWIDTH'b1111111001101110,
        `W_DATA_BITWIDTH'b0000000101011110,
        `W_DATA_BITWIDTH'b1111111011001011,
        `W_DATA_BITWIDTH'b0000001101111000,
        `W_DATA_BITWIDTH'b0000011010000001,
        `W_DATA_BITWIDTH'b1111100010110110,
        `W_DATA_BITWIDTH'b1111110111010110,
        `W_DATA_BITWIDTH'b0000011010111110,
        `W_DATA_BITWIDTH'b1111101110100010,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b0000001000000110,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111100010100101,
        `W_DATA_BITWIDTH'b1111111011100000,
        `W_DATA_BITWIDTH'b0000001110100010,
        `W_DATA_BITWIDTH'b0000000111011111,
        `W_DATA_BITWIDTH'b1111110010111011,
        `W_DATA_BITWIDTH'b0000010000100101,
        `W_DATA_BITWIDTH'b0000010000100101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_DATA_BITWIDTH'b1111111101010101,
        `W_DATA_BITWIDTH'b0000000011101111,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110101011010,
        `W_DATA_BITWIDTH'b1111110101010100,
        `W_DATA_BITWIDTH'b0000001011110011,
        `W_DATA_BITWIDTH'b1111111001100101,
        `W_DATA_BITWIDTH'b0000010101111110,
        `W_DATA_BITWIDTH'b0000010010100101,
        `W_DATA_BITWIDTH'b1111011110010000,
        `W_DATA_BITWIDTH'b1111110001000001,
        `W_DATA_BITWIDTH'b0000001101001011,
        `W_DATA_BITWIDTH'b0000011001011010,
        `W_DATA_BITWIDTH'b1111100001111110,
        `W_DATA_BITWIDTH'b0000010010100111,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b1111111000111101,
        `W_DATA_BITWIDTH'b1111111011111100,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000110001000,
        `W_DATA_BITWIDTH'b1111110011001010,
        `W_DATA_BITWIDTH'b1111111001000011,
        `W_DATA_BITWIDTH'b1111111001011001,
        `W_DATA_BITWIDTH'b0000001010000101,
        `W_DATA_BITWIDTH'b0000001100001100,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111111001001011,
        `W_DATA_BITWIDTH'b0000010001001101,
        `W_DATA_BITWIDTH'b0000100000011111,
        `W_DATA_BITWIDTH'b1111100000100000,
        `W_DATA_BITWIDTH'b1111100111110111,
        `W_DATA_BITWIDTH'b0000001011100001,
        `W_DATA_BITWIDTH'b1111111101101011,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b0000001010100100,
        `W_DATA_BITWIDTH'b1111111000111110,
        `W_DATA_BITWIDTH'b0000001000000011,
        `W_DATA_BITWIDTH'b1111110101011011,
        `W_DATA_BITWIDTH'b1111111011010100,
        `W_DATA_BITWIDTH'b0000010010110001,
        `W_DATA_BITWIDTH'b1111110110001010,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b0000001110100101,
        `W_DATA_BITWIDTH'b0000000011100100,
        `W_DATA_BITWIDTH'b0000000111101001,
        `W_DATA_BITWIDTH'b0000001110011000,
        `W_DATA_BITWIDTH'b1111111101101010,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000001100101010,
        `W_DATA_BITWIDTH'b0000001001011111,
        `W_DATA_BITWIDTH'b1111111001010011,
        `W_DATA_BITWIDTH'b1111101010010111,
        `W_DATA_BITWIDTH'b1111110010010011,
        `W_DATA_BITWIDTH'b0000001111110100,
        `W_DATA_BITWIDTH'b0000000111011011,
        `W_DATA_BITWIDTH'b0000001011110101,
        `W_DATA_BITWIDTH'b1111100111101101,
        `W_DATA_BITWIDTH'b0000100000011000,
        `W_DATA_BITWIDTH'b1111111011111101,
        `W_DATA_BITWIDTH'b1111111011111101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_DATA_BITWIDTH'b1111110101111111,
        `W_DATA_BITWIDTH'b1111111001010010,
        `W_DATA_BITWIDTH'b1111110101000101,
        `W_DATA_BITWIDTH'b0000000110011101,
        `W_DATA_BITWIDTH'b1111111100000001,
        `W_DATA_BITWIDTH'b0000001110111001,
        `W_DATA_BITWIDTH'b0000001100010101,
        `W_DATA_BITWIDTH'b1111111000101001,
        `W_DATA_BITWIDTH'b1111110001010101,
        `W_DATA_BITWIDTH'b1111110110000011,
        `W_DATA_BITWIDTH'b1111111010110011,
        `W_DATA_BITWIDTH'b1111110000110011,
        `W_DATA_BITWIDTH'b1111110011010001,
        `W_DATA_BITWIDTH'b0000001110101010,
        `W_DATA_BITWIDTH'b0000010000011111,
        `W_DATA_BITWIDTH'b1111111010011010,
        `W_DATA_BITWIDTH'b0000000110010000,
        `W_DATA_BITWIDTH'b1111110100011101,
        `W_DATA_BITWIDTH'b0000001010011111,
        `W_DATA_BITWIDTH'b1111111000000011,
        `W_DATA_BITWIDTH'b1111111000111100,
        `W_DATA_BITWIDTH'b1111111011010000,
        `W_DATA_BITWIDTH'b0000001011001111,
        `W_DATA_BITWIDTH'b1111110110100001,
        `W_DATA_BITWIDTH'b1111101011111100,
        `W_DATA_BITWIDTH'b1111110110101110,
        `W_DATA_BITWIDTH'b0000001110000011,
        `W_DATA_BITWIDTH'b1111111100000101,
        `W_DATA_BITWIDTH'b0000000101110010,
        `W_DATA_BITWIDTH'b1111110000011010,
        `W_DATA_BITWIDTH'b0000000101011101,
        `W_DATA_BITWIDTH'b1111111001101101,
        `W_DATA_BITWIDTH'b0000001101101101,
        `W_DATA_BITWIDTH'b1111110101111010,
        `W_DATA_BITWIDTH'b0000000100000000,
        `W_DATA_BITWIDTH'b1111111010111101,
        `W_DATA_BITWIDTH'b1111110010101100,
        `W_DATA_BITWIDTH'b0000001011111000,
        `W_DATA_BITWIDTH'b1111110011100100,
        `W_DATA_BITWIDTH'b1111110100001011,
        `W_DATA_BITWIDTH'b1111110110001100,
        `W_DATA_BITWIDTH'b1111100111101010,
        `W_DATA_BITWIDTH'b1111110101001111,
        `W_DATA_BITWIDTH'b1111111011011010,
        `W_DATA_BITWIDTH'b1111111000101110,
        `W_DATA_BITWIDTH'b0000000110100011,
        `W_DATA_BITWIDTH'b1111110011011100,
        `W_DATA_BITWIDTH'b1111110011010001,
        `W_DATA_BITWIDTH'b1111110111000100,
        `W_DATA_BITWIDTH'b0000001100001101,
        `W_DATA_BITWIDTH'b1111111001110101,
        `W_DATA_BITWIDTH'b1111110111000100,
        `W_DATA_BITWIDTH'b0000001100010111,
        `W_DATA_BITWIDTH'b1111111000000011,
        `W_DATA_BITWIDTH'b1111110000101111,
        `W_DATA_BITWIDTH'b1111100110110000,
        `W_DATA_BITWIDTH'b0000010111000111,
        `W_DATA_BITWIDTH'b1111110111111101,
        `W_DATA_BITWIDTH'b0000001100100010,
        `W_DATA_BITWIDTH'b1111110111101110,
        `W_DATA_BITWIDTH'b1111111010111101,
        `W_DATA_BITWIDTH'b1111111011000010,
        `W_DATA_BITWIDTH'b1111110001100110,
        `W_DATA_BITWIDTH'b0000001000110111,
        `W_DATA_BITWIDTH'b1111110011000011,
        `W_DATA_BITWIDTH'b0000000111100000,
        `W_DATA_BITWIDTH'b1111101111011111,
        `W_DATA_BITWIDTH'b1111101000111111,
        `W_DATA_BITWIDTH'b0000001011010011,
        `W_DATA_BITWIDTH'b1111111001110100,
        `W_DATA_BITWIDTH'b0000001010011001,
        `W_DATA_BITWIDTH'b1111110011100111,
        `W_DATA_BITWIDTH'b0000001011011111,
        `W_DATA_BITWIDTH'b1111110110000101,
        `W_DATA_BITWIDTH'b1111110111010100,
        `W_DATA_BITWIDTH'b0000010100001001,
        `W_DATA_BITWIDTH'b1111110110100100,
        `W_DATA_BITWIDTH'b0000010000011101,
        `W_DATA_BITWIDTH'b0000001010111011,
        `W_DATA_BITWIDTH'b0000001000001010,
        `W_DATA_BITWIDTH'b0000000111000000,
        `W_DATA_BITWIDTH'b0000000110000101,
        `W_DATA_BITWIDTH'b1111100111110100,
        `W_DATA_BITWIDTH'b1111101010010100,
        `W_DATA_BITWIDTH'b0000010001010101,
        `W_DATA_BITWIDTH'b0000000110100000,
        `W_DATA_BITWIDTH'b1111111011011011,
        `W_DATA_BITWIDTH'b1111110110100100,
        `W_DATA_BITWIDTH'b1111101000100111,
        `W_DATA_BITWIDTH'b0000000101101101,
        `W_DATA_BITWIDTH'b0000001000010000,
        `W_DATA_BITWIDTH'b0000010100010001,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b0000001100110110,
        `W_DATA_BITWIDTH'b0000000110000001,
        `W_DATA_BITWIDTH'b0000010010110000,
        `W_DATA_BITWIDTH'b1111110001100110,
        `W_DATA_BITWIDTH'b0000000101011011,
        `W_DATA_BITWIDTH'b0000001100101000,
        `W_DATA_BITWIDTH'b1111110001011011,
        `W_DATA_BITWIDTH'b1111111000011101,
        `W_DATA_BITWIDTH'b0000001011010001,
        `W_DATA_BITWIDTH'b0000011000001010,
        `W_DATA_BITWIDTH'b1111110011001011,
        `W_DATA_BITWIDTH'b1111111000000001,
        `W_DATA_BITWIDTH'b1111110111100001,
        `W_DATA_BITWIDTH'b1111110100111000,
        `W_DATA_BITWIDTH'b0000000101010000,
        `W_DATA_BITWIDTH'b0000000111111000,
        `W_DATA_BITWIDTH'b1111110011101100,
        `W_DATA_BITWIDTH'b1111110110110100,
        `W_DATA_BITWIDTH'b0000001100001000,
        `W_DATA_BITWIDTH'b0000001101111010,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b0000000101110101,
        `W_DATA_BITWIDTH'b0000000101001110,
        `W_DATA_BITWIDTH'b0000000100111010,
        `W_DATA_BITWIDTH'b0000001100011100,
        `W_DATA_BITWIDTH'b1111111010010010,
        `W_DATA_BITWIDTH'b0000000011111110,
        `W_DATA_BITWIDTH'b1111110100000011,
        `W_DATA_BITWIDTH'b1111110101111100,
        `W_DATA_BITWIDTH'b1111101111101010,
        `W_DATA_BITWIDTH'b1111101100111011,
        `W_DATA_BITWIDTH'b1111110011100110,
        `W_DATA_BITWIDTH'b1111101010110101,
        `W_DATA_BITWIDTH'b1111101100110010,
        `W_DATA_BITWIDTH'b1111111000000011,
        `W_DATA_BITWIDTH'b1111111010010111,
        `W_DATA_BITWIDTH'b0000000101011100,
        `W_DATA_BITWIDTH'b0000000101011100
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_DATA_BITWIDTH'b0000000101000011,
        `W_DATA_BITWIDTH'b0000001101011111,
        `W_DATA_BITWIDTH'b0000010111001011,
        `W_DATA_BITWIDTH'b0000001111100110,
        `W_DATA_BITWIDTH'b0000010000111011,
        `W_DATA_BITWIDTH'b0000000111111111,
        `W_DATA_BITWIDTH'b0000001110001001,
        `W_DATA_BITWIDTH'b1111111001010100,
        `W_DATA_BITWIDTH'b1111111010100001,
        `W_DATA_BITWIDTH'b1111101110111101,
        `W_DATA_BITWIDTH'b1111101010110101,
        `W_DATA_BITWIDTH'b1111101110000011,
        `W_DATA_BITWIDTH'b1111110111111100,
        `W_DATA_BITWIDTH'b1111110110000011,
        `W_DATA_BITWIDTH'b1111110100110101,
        `W_DATA_BITWIDTH'b1111110101011001,
        `W_DATA_BITWIDTH'b0000001111001011,
        `W_DATA_BITWIDTH'b0000000110011100,
        `W_DATA_BITWIDTH'b1111111011100001,
        `W_DATA_BITWIDTH'b1111110110100111,
        `W_DATA_BITWIDTH'b0000001000110101,
        `W_DATA_BITWIDTH'b1111110100101010,
        `W_DATA_BITWIDTH'b1111110010100000,
        `W_DATA_BITWIDTH'b1111101111100000,
        `W_DATA_BITWIDTH'b0000000100001111,
        `W_DATA_BITWIDTH'b0000000111110001,
        `W_DATA_BITWIDTH'b0000000111111010,
        `W_DATA_BITWIDTH'b0000010010100100,
        `W_DATA_BITWIDTH'b0000001101101100,
        `W_DATA_BITWIDTH'b0000001001011011,
        `W_DATA_BITWIDTH'b1111110101011110,
        `W_DATA_BITWIDTH'b1111110010110001,
        `W_DATA_BITWIDTH'b0000001000111001,
        `W_DATA_BITWIDTH'b0000000110000001,
        `W_DATA_BITWIDTH'b1111101111101101,
        `W_DATA_BITWIDTH'b0000001100100001,
        `W_DATA_BITWIDTH'b0000001111001011,
        `W_DATA_BITWIDTH'b0000001011000110,
        `W_DATA_BITWIDTH'b1111101101011101,
        `W_DATA_BITWIDTH'b0000001010010011,
        `W_DATA_BITWIDTH'b1111111011111001,
        `W_DATA_BITWIDTH'b1111111010110101,
        `W_DATA_BITWIDTH'b1111111000011111,
        `W_DATA_BITWIDTH'b1111111011010100,
        `W_DATA_BITWIDTH'b1111110000000000,
        `W_DATA_BITWIDTH'b0000001001111100,
        `W_DATA_BITWIDTH'b0000001000010101,
        `W_DATA_BITWIDTH'b0000001011010101,
        `W_DATA_BITWIDTH'b1111110011111011,
        `W_DATA_BITWIDTH'b1111101110011001,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b0000000101011110,
        `W_DATA_BITWIDTH'b1111110110001000,
        `W_DATA_BITWIDTH'b0000001000111101,
        `W_DATA_BITWIDTH'b1111110110111111,
        `W_DATA_BITWIDTH'b0000000111101001,
        `W_DATA_BITWIDTH'b0000001001011001,
        `W_DATA_BITWIDTH'b1111110111111101,
        `W_DATA_BITWIDTH'b0000001010101100,
        `W_DATA_BITWIDTH'b0000000101000001,
        `W_DATA_BITWIDTH'b1111110010110101,
        `W_DATA_BITWIDTH'b1111110111001011,
        `W_DATA_BITWIDTH'b1111111000111101,
        `W_DATA_BITWIDTH'b0000001000110100,
        `W_DATA_BITWIDTH'b1111111000110000,
        `W_DATA_BITWIDTH'b0000000100111010,
        `W_DATA_BITWIDTH'b1111111011011101,
        `W_DATA_BITWIDTH'b0000001000111100,
        `W_DATA_BITWIDTH'b1111111000100011,
        `W_DATA_BITWIDTH'b0000001000111000,
        `W_DATA_BITWIDTH'b1111110100100010,
        `W_DATA_BITWIDTH'b1111110001110100,
        `W_DATA_BITWIDTH'b1111101101011011,
        `W_DATA_BITWIDTH'b1111110101100010,
        `W_DATA_BITWIDTH'b1111110101101110,
        `W_DATA_BITWIDTH'b1111111001010100,
        `W_DATA_BITWIDTH'b1111110101100101,
        `W_DATA_BITWIDTH'b0000000110110111,
        `W_DATA_BITWIDTH'b0000001001111101,
        `W_DATA_BITWIDTH'b1111111000011100,
        `W_DATA_BITWIDTH'b0000000101010011,
        `W_DATA_BITWIDTH'b1111110100001100,
        `W_DATA_BITWIDTH'b0000010000011100,
        `W_DATA_BITWIDTH'b1111110101111001,
        `W_DATA_BITWIDTH'b0000000101000101,
        `W_DATA_BITWIDTH'b0000000111101011,
        `W_DATA_BITWIDTH'b1111110111000111,
        `W_DATA_BITWIDTH'b1111111000111100,
        `W_DATA_BITWIDTH'b0000001101100011,
        `W_DATA_BITWIDTH'b1111110101010010,
        `W_DATA_BITWIDTH'b1111110110101111,
        `W_DATA_BITWIDTH'b0000000101011010,
        `W_DATA_BITWIDTH'b0000000100110100,
        `W_DATA_BITWIDTH'b1111110101100110,
        `W_DATA_BITWIDTH'b1111111100000011,
        `W_DATA_BITWIDTH'b0000000111110001,
        `W_DATA_BITWIDTH'b1111111011111111,
        `W_DATA_BITWIDTH'b1111110101100111,
        `W_DATA_BITWIDTH'b0000001100101110,
        `W_DATA_BITWIDTH'b0000000110011011,
        `W_DATA_BITWIDTH'b0000001011100111,
        `W_DATA_BITWIDTH'b1111110010110011,
        `W_DATA_BITWIDTH'b0000010101110101,
        `W_DATA_BITWIDTH'b0000001001011111,
        `W_DATA_BITWIDTH'b0000000100010111,
        `W_DATA_BITWIDTH'b1111100101101101,
        `W_DATA_BITWIDTH'b1111110100010010,
        `W_DATA_BITWIDTH'b0000001110100000,
        `W_DATA_BITWIDTH'b1111110011101110,
        `W_DATA_BITWIDTH'b0000000100110111,
        `W_DATA_BITWIDTH'b1111110010110100,
        `W_DATA_BITWIDTH'b0000000100010100,
        `W_DATA_BITWIDTH'b1111101111110101,
        `W_DATA_BITWIDTH'b1111111011011011,
        `W_DATA_BITWIDTH'b1111101010010001,
        `W_DATA_BITWIDTH'b0000010010001110,
        `W_DATA_BITWIDTH'b0000001101011111,
        `W_DATA_BITWIDTH'b1111101000100110,
        `W_DATA_BITWIDTH'b1111110101010111,
        `W_DATA_BITWIDTH'b0000001001010010,
        `W_DATA_BITWIDTH'b0000001001111010,
        `W_DATA_BITWIDTH'b1111110101110001,
        `W_DATA_BITWIDTH'b0000001000011000,
        `W_DATA_BITWIDTH'b0000001111011011,
        `W_DATA_BITWIDTH'b0000001111011011,
        `W_DATA_BITWIDTH'b0000001101101001,
        `W_DATA_BITWIDTH'b0000010010001000,
        `W_DATA_BITWIDTH'b0000001010011001,
        `W_DATA_BITWIDTH'b0000001011000011,
        `W_DATA_BITWIDTH'b0000001100001010,
        `W_DATA_BITWIDTH'b1111110100110010,
        `W_DATA_BITWIDTH'b1111111001111000,
        `W_DATA_BITWIDTH'b1111110100110100,
        `W_DATA_BITWIDTH'b1111111010101110,
        `W_DATA_BITWIDTH'b1111111000011000,
        `W_DATA_BITWIDTH'b0000001000101100,
        `W_DATA_BITWIDTH'b1111110100101100,
        `W_DATA_BITWIDTH'b1111110100100111,
        `W_DATA_BITWIDTH'b0000001100010010,
        `W_DATA_BITWIDTH'b1111111010111110,
        `W_DATA_BITWIDTH'b1111111010111110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_DATA_BITWIDTH'b1111110101111000,
        `W_DATA_BITWIDTH'b0000001100011110,
        `W_DATA_BITWIDTH'b0000001111111111,
        `W_DATA_BITWIDTH'b1111110011111001,
        `W_DATA_BITWIDTH'b1111110110000100,
        `W_DATA_BITWIDTH'b0000000111111100,
        `W_DATA_BITWIDTH'b1111101111000110,
        `W_DATA_BITWIDTH'b1111110110010110,
        `W_DATA_BITWIDTH'b1111110000101110,
        `W_DATA_BITWIDTH'b0000010001010110,
        `W_DATA_BITWIDTH'b1111101010001110,
        `W_DATA_BITWIDTH'b1111111011110011,
        `W_DATA_BITWIDTH'b0000001000110001,
        `W_DATA_BITWIDTH'b1111111011001100,
        `W_DATA_BITWIDTH'b0000010000001111,
        `W_DATA_BITWIDTH'b1111101111100111,
        `W_DATA_BITWIDTH'b0000001000111011,
        `W_DATA_BITWIDTH'b1111111000001010,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b1111111011111010,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b1111110101011011,
        `W_DATA_BITWIDTH'b1111110011100001,
        `W_DATA_BITWIDTH'b1111110011010111,
        `W_DATA_BITWIDTH'b1111110001101011,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b1111110000101010,
        `W_DATA_BITWIDTH'b1111110101010010,
        `W_DATA_BITWIDTH'b1111111010000111,
        `W_DATA_BITWIDTH'b0000010001000110,
        `W_DATA_BITWIDTH'b0000000101010101,
        `W_DATA_BITWIDTH'b0000000011111110,
        `W_DATA_BITWIDTH'b0000000100011010,
        `W_DATA_BITWIDTH'b1111111000111001,
        `W_DATA_BITWIDTH'b0000000100011111,
        `W_DATA_BITWIDTH'b1111101111001110,
        `W_DATA_BITWIDTH'b0000000100101001,
        `W_DATA_BITWIDTH'b0000001011110001,
        `W_DATA_BITWIDTH'b0000001100011001,
        `W_DATA_BITWIDTH'b0000000100100100,
        `W_DATA_BITWIDTH'b1111110011000110,
        `W_DATA_BITWIDTH'b0000000111010110,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b0000010000000100,
        `W_DATA_BITWIDTH'b0000000101000010,
        `W_DATA_BITWIDTH'b1111111010000110,
        `W_DATA_BITWIDTH'b1111111010110111,
        `W_DATA_BITWIDTH'b0000000110011010,
        `W_DATA_BITWIDTH'b1111110101001100,
        `W_DATA_BITWIDTH'b1111110111000010,
        `W_DATA_BITWIDTH'b1111111010110011,
        `W_DATA_BITWIDTH'b1111111001101110,
        `W_DATA_BITWIDTH'b0000001110110101,
        `W_DATA_BITWIDTH'b1111111001111011,
        `W_DATA_BITWIDTH'b0000000101000001,
        `W_DATA_BITWIDTH'b0000000101010111,
        `W_DATA_BITWIDTH'b1111110111101111,
        `W_DATA_BITWIDTH'b1111101110001100,
        `W_DATA_BITWIDTH'b1111110010000111,
        `W_DATA_BITWIDTH'b0000001010111010,
        `W_DATA_BITWIDTH'b0000001000110110,
        `W_DATA_BITWIDTH'b1111110100110110,
        `W_DATA_BITWIDTH'b1111110000110010,
        `W_DATA_BITWIDTH'b1111111010100001,
        `W_DATA_BITWIDTH'b1111110011101110,
        `W_DATA_BITWIDTH'b1111110111100101,
        `W_DATA_BITWIDTH'b1111111001101101,
        `W_DATA_BITWIDTH'b1111101101101000,
        `W_DATA_BITWIDTH'b0000001000100110,
        `W_DATA_BITWIDTH'b1111110011110101,
        `W_DATA_BITWIDTH'b0000010100111111,
        `W_DATA_BITWIDTH'b0000000101110111,
        `W_DATA_BITWIDTH'b1111101111101011,
        `W_DATA_BITWIDTH'b1111110001001100,
        `W_DATA_BITWIDTH'b0000011010110011,
        `W_DATA_BITWIDTH'b1111111011010101,
        `W_DATA_BITWIDTH'b0000010011111011,
        `W_DATA_BITWIDTH'b1111111001011110,
        `W_DATA_BITWIDTH'b0000000100001010,
        `W_DATA_BITWIDTH'b1111111010111100,
        `W_DATA_BITWIDTH'b0000001100010001,
        `W_DATA_BITWIDTH'b0000011011000000,
        `W_DATA_BITWIDTH'b1111111000010000,
        `W_DATA_BITWIDTH'b0000000100011101,
        `W_DATA_BITWIDTH'b1111110111100001,
        `W_DATA_BITWIDTH'b1111101001110000,
        `W_DATA_BITWIDTH'b1111110110011111,
        `W_DATA_BITWIDTH'b1111110000101010,
        `W_DATA_BITWIDTH'b0000000101000101,
        `W_DATA_BITWIDTH'b0000001000100001,
        `W_DATA_BITWIDTH'b0000000101110000,
        `W_DATA_BITWIDTH'b1111110011110011,
        `W_DATA_BITWIDTH'b0000001010111101,
        `W_DATA_BITWIDTH'b1111111011000101,
        `W_DATA_BITWIDTH'b1111111011100010,
        `W_DATA_BITWIDTH'b1111111010111100,
        `W_DATA_BITWIDTH'b1111111010001000,
        `W_DATA_BITWIDTH'b1111110111110000,
        `W_DATA_BITWIDTH'b0000000100011111,
        `W_DATA_BITWIDTH'b1111111001001000,
        `W_DATA_BITWIDTH'b0000000101011100,
        `W_DATA_BITWIDTH'b1111100100101101,
        `W_DATA_BITWIDTH'b1111110111001101,
        `W_DATA_BITWIDTH'b1111110100001110,
        `W_DATA_BITWIDTH'b1111111001000000,
        `W_DATA_BITWIDTH'b0000000100000011,
        `W_DATA_BITWIDTH'b1111110110111111,
        `W_DATA_BITWIDTH'b1111101000010110,
        `W_DATA_BITWIDTH'b0000001000001011,
        `W_DATA_BITWIDTH'b0000010001011111,
        `W_DATA_BITWIDTH'b1111110111001010,
        `W_DATA_BITWIDTH'b1111110010101101,
        `W_DATA_BITWIDTH'b0000010010101011,
        `W_DATA_BITWIDTH'b0000001001100111,
        `W_DATA_BITWIDTH'b1111111000011001,
        `W_DATA_BITWIDTH'b1111101011111101,
        `W_DATA_BITWIDTH'b1111110110100010,
        `W_DATA_BITWIDTH'b1111111000000110,
        `W_DATA_BITWIDTH'b0000001001000101,
        `W_DATA_BITWIDTH'b1111111011110010,
        `W_DATA_BITWIDTH'b0000000100001001,
        `W_DATA_BITWIDTH'b0000000100111110,
        `W_DATA_BITWIDTH'b1111110111110000,
        `W_DATA_BITWIDTH'b1111110100101101,
        `W_DATA_BITWIDTH'b0000000101001111,
        `W_DATA_BITWIDTH'b0000001001001011,
        `W_DATA_BITWIDTH'b1111110010001011,
        `W_DATA_BITWIDTH'b1111110010110111,
        `W_DATA_BITWIDTH'b1111111011111010,
        `W_DATA_BITWIDTH'b1111111011100000,
        `W_DATA_BITWIDTH'b1111111011100000
    };

// w_c_idx
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00110
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00110
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00110
    };

// w_r_idx
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };

// w_k_idx
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };

// w_pos_ptr
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000011,
        `W_POS_PTR_BITWIDTH'b00000000110,
        `W_POS_PTR_BITWIDTH'b00000001001,
        `W_POS_PTR_BITWIDTH'b00000001100,
        `W_POS_PTR_BITWIDTH'b00000001111,
        `W_POS_PTR_BITWIDTH'b00000010010,
        `W_POS_PTR_BITWIDTH'b00000010101,
        `W_POS_PTR_BITWIDTH'b00000011000,
        `W_POS_PTR_BITWIDTH'b00000011011,
        `W_POS_PTR_BITWIDTH'b00000011110,
        `W_POS_PTR_BITWIDTH'b00000100001,
        `W_POS_PTR_BITWIDTH'b00000100100,
        `W_POS_PTR_BITWIDTH'b00000100110,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000101010,
        `W_POS_PTR_BITWIDTH'b00000101101,
        `W_POS_PTR_BITWIDTH'b00000110000,
        `W_POS_PTR_BITWIDTH'b00000110011,
        `W_POS_PTR_BITWIDTH'b00000110110,
        `W_POS_PTR_BITWIDTH'b00000111001,
        `W_POS_PTR_BITWIDTH'b00000111011,
        `W_POS_PTR_BITWIDTH'b00000111110,
        `W_POS_PTR_BITWIDTH'b00000111110
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00001000100,
        `W_POS_PTR_BITWIDTH'b00001000111,
        `W_POS_PTR_BITWIDTH'b00001001001,
        `W_POS_PTR_BITWIDTH'b00001001100,
        `W_POS_PTR_BITWIDTH'b00001001111,
        `W_POS_PTR_BITWIDTH'b00001010001,
        `W_POS_PTR_BITWIDTH'b00001010100,
        `W_POS_PTR_BITWIDTH'b00001010111,
        `W_POS_PTR_BITWIDTH'b00001011000,
        `W_POS_PTR_BITWIDTH'b00001011011,
        `W_POS_PTR_BITWIDTH'b00001011110,
        `W_POS_PTR_BITWIDTH'b00001100001,
        `W_POS_PTR_BITWIDTH'b00001100100,
        `W_POS_PTR_BITWIDTH'b00001100111,
        `W_POS_PTR_BITWIDTH'b00001101010,
        `W_POS_PTR_BITWIDTH'b00001101101,
        `W_POS_PTR_BITWIDTH'b00001110000,
        `W_POS_PTR_BITWIDTH'b00001110011,
        `W_POS_PTR_BITWIDTH'b00001110110,
        `W_POS_PTR_BITWIDTH'b00001111001,
        `W_POS_PTR_BITWIDTH'b00001111100,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010000010,
        `W_POS_PTR_BITWIDTH'b00010000010
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00010000110,
        `W_POS_PTR_BITWIDTH'b00010001001,
        `W_POS_PTR_BITWIDTH'b00010001010,
        `W_POS_PTR_BITWIDTH'b00010001100,
        `W_POS_PTR_BITWIDTH'b00010001111,
        `W_POS_PTR_BITWIDTH'b00010010001,
        `W_POS_PTR_BITWIDTH'b00010010100,
        `W_POS_PTR_BITWIDTH'b00010010111,
        `W_POS_PTR_BITWIDTH'b00010011010,
        `W_POS_PTR_BITWIDTH'b00010011100,
        `W_POS_PTR_BITWIDTH'b00010011111,
        `W_POS_PTR_BITWIDTH'b00010100010,
        `W_POS_PTR_BITWIDTH'b00010100101,
        `W_POS_PTR_BITWIDTH'b00010100110,
        `W_POS_PTR_BITWIDTH'b00010101000,
        `W_POS_PTR_BITWIDTH'b00010101001,
        `W_POS_PTR_BITWIDTH'b00010101100,
        `W_POS_PTR_BITWIDTH'b00010101111,
        `W_POS_PTR_BITWIDTH'b00010110010,
        `W_POS_PTR_BITWIDTH'b00010110101,
        `W_POS_PTR_BITWIDTH'b00010110110,
        `W_POS_PTR_BITWIDTH'b00010111001,
        `W_POS_PTR_BITWIDTH'b00010111100,
        `W_POS_PTR_BITWIDTH'b00010111100
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000101,
        `W_POS_PTR_BITWIDTH'b00000001011,
        `W_POS_PTR_BITWIDTH'b00000010000,
        `W_POS_PTR_BITWIDTH'b00000010110,
        `W_POS_PTR_BITWIDTH'b00000011010,
        `W_POS_PTR_BITWIDTH'b00000100001,
        `W_POS_PTR_BITWIDTH'b00000100010,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000101111,
        `W_POS_PTR_BITWIDTH'b00000110011,
        `W_POS_PTR_BITWIDTH'b00000110111,
        `W_POS_PTR_BITWIDTH'b00000111101,
        `W_POS_PTR_BITWIDTH'b00001000010,
        `W_POS_PTR_BITWIDTH'b00001001000,
        `W_POS_PTR_BITWIDTH'b00001001110,
        `W_POS_PTR_BITWIDTH'b00001010101,
        `W_POS_PTR_BITWIDTH'b00001011010,
        `W_POS_PTR_BITWIDTH'b00001011101,
        `W_POS_PTR_BITWIDTH'b00001100100,
        `W_POS_PTR_BITWIDTH'b00001101010,
        `W_POS_PTR_BITWIDTH'b00001101111,
        `W_POS_PTR_BITWIDTH'b00001110101,
        `W_POS_PTR_BITWIDTH'b00001110101
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00010000011,
        `W_POS_PTR_BITWIDTH'b00010001010,
        `W_POS_PTR_BITWIDTH'b00010010010,
        `W_POS_PTR_BITWIDTH'b00010010101,
        `W_POS_PTR_BITWIDTH'b00010011010,
        `W_POS_PTR_BITWIDTH'b00010011111,
        `W_POS_PTR_BITWIDTH'b00010100010,
        `W_POS_PTR_BITWIDTH'b00010101000,
        `W_POS_PTR_BITWIDTH'b00010110000,
        `W_POS_PTR_BITWIDTH'b00010110110,
        `W_POS_PTR_BITWIDTH'b00010111010,
        `W_POS_PTR_BITWIDTH'b00011000000,
        `W_POS_PTR_BITWIDTH'b00011000110,
        `W_POS_PTR_BITWIDTH'b00011001101,
        `W_POS_PTR_BITWIDTH'b00011010101,
        `W_POS_PTR_BITWIDTH'b00011011001,
        `W_POS_PTR_BITWIDTH'b00011011111,
        `W_POS_PTR_BITWIDTH'b00011100100,
        `W_POS_PTR_BITWIDTH'b00011101100,
        `W_POS_PTR_BITWIDTH'b00011110010,
        `W_POS_PTR_BITWIDTH'b00011111000,
        `W_POS_PTR_BITWIDTH'b00011111101,
        `W_POS_PTR_BITWIDTH'b00100000011,
        `W_POS_PTR_BITWIDTH'b00100000011
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00100010000,
        `W_POS_PTR_BITWIDTH'b00100010101,
        `W_POS_PTR_BITWIDTH'b00100011100,
        `W_POS_PTR_BITWIDTH'b00100100010,
        `W_POS_PTR_BITWIDTH'b00100100110,
        `W_POS_PTR_BITWIDTH'b00100101011,
        `W_POS_PTR_BITWIDTH'b00100101111,
        `W_POS_PTR_BITWIDTH'b00100110111,
        `W_POS_PTR_BITWIDTH'b00100111101,
        `W_POS_PTR_BITWIDTH'b00101000011,
        `W_POS_PTR_BITWIDTH'b00101001001,
        `W_POS_PTR_BITWIDTH'b00101001111,
        `W_POS_PTR_BITWIDTH'b00101010101,
        `W_POS_PTR_BITWIDTH'b00101011100,
        `W_POS_PTR_BITWIDTH'b00101100001,
        `W_POS_PTR_BITWIDTH'b00101100110,
        `W_POS_PTR_BITWIDTH'b00101101100,
        `W_POS_PTR_BITWIDTH'b00101101111,
        `W_POS_PTR_BITWIDTH'b00101110100,
        `W_POS_PTR_BITWIDTH'b00101111011,
        `W_POS_PTR_BITWIDTH'b00110000000,
        `W_POS_PTR_BITWIDTH'b00110000101,
        `W_POS_PTR_BITWIDTH'b00110001000,
        `W_POS_PTR_BITWIDTH'b00110001000
    };

// w_all
