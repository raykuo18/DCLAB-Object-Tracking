// w_c_idx
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00101
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00011,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00110,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00100,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00101,
        `W_C_BITWIDTH'b00111,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };

// w_c_idx
