// w_data
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_DATA_BITWIDTH'b1111110011100101,
        `W_DATA_BITWIDTH'b1111111001011110,
        `W_DATA_BITWIDTH'b0000001001011101,
        `W_DATA_BITWIDTH'b1111111101011000,
        `W_DATA_BITWIDTH'b1111110101101101,
        `W_DATA_BITWIDTH'b1111110010110110,
        `W_DATA_BITWIDTH'b0000001110111010,
        `W_DATA_BITWIDTH'b1111111010001100,
        `W_DATA_BITWIDTH'b0000001000001011,
        `W_DATA_BITWIDTH'b1111101111110111,
        `W_DATA_BITWIDTH'b0000000010111010,
        `W_DATA_BITWIDTH'b0000001101011100,
        `W_DATA_BITWIDTH'b0000000110001011,
        `W_DATA_BITWIDTH'b1111110000101100,
        `W_DATA_BITWIDTH'b0000001110000100,
        `W_DATA_BITWIDTH'b0000010011010001,
        `W_DATA_BITWIDTH'b1111100001100110,
        `W_DATA_BITWIDTH'b0000001110000111,
        `W_DATA_BITWIDTH'b1111110110101001,
        `W_DATA_BITWIDTH'b1111111000011000,
        `W_DATA_BITWIDTH'b0000001000010001,
        `W_DATA_BITWIDTH'b0000000110110111,
        `W_DATA_BITWIDTH'b0000000010000000,
        `W_DATA_BITWIDTH'b1111110100000000,
        `W_DATA_BITWIDTH'b0000000110010101,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b0000000101011011,
        `W_DATA_BITWIDTH'b0000001000101100,
        `W_DATA_BITWIDTH'b0000000111010100,
        `W_DATA_BITWIDTH'b1111111000001000,
        `W_DATA_BITWIDTH'b1111111011011010,
        `W_DATA_BITWIDTH'b0000000010011110,
        `W_DATA_BITWIDTH'b1111111100110001,
        `W_DATA_BITWIDTH'b0000010000101111,
        `W_DATA_BITWIDTH'b1111101001000011,
        `W_DATA_BITWIDTH'b1111111000011101,
        `W_DATA_BITWIDTH'b1111110010111111,
        `W_DATA_BITWIDTH'b1111111101110010,
        `W_DATA_BITWIDTH'b1111111011110001,
        `W_DATA_BITWIDTH'b1111111011100011,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000111100110,
        `W_DATA_BITWIDTH'b0000010001100000,
        `W_DATA_BITWIDTH'b1111101101100010,
        `W_DATA_BITWIDTH'b1111111101110110,
        `W_DATA_BITWIDTH'b0000001110000101,
        `W_DATA_BITWIDTH'b1111100111001110,
        `W_DATA_BITWIDTH'b0000000101011000,
        `W_DATA_BITWIDTH'b0000001101011101,
        `W_DATA_BITWIDTH'b1111110000000010,
        `W_DATA_BITWIDTH'b0000001000001000,
        `W_DATA_BITWIDTH'b1111100111110100,
        `W_DATA_BITWIDTH'b0000000111100011,
        `W_DATA_BITWIDTH'b0000001001010101,
        `W_DATA_BITWIDTH'b0000000100011010,
        `W_DATA_BITWIDTH'b0000010011000111,
        `W_DATA_BITWIDTH'b0000000010000001,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000000011100001,
        `W_DATA_BITWIDTH'b1111111010100101,
        `W_DATA_BITWIDTH'b0000000101001001,
        `W_DATA_BITWIDTH'b0000001111100110,
        `W_DATA_BITWIDTH'b0000001010101001,
        `W_DATA_BITWIDTH'b0000011011010011,
        `W_DATA_BITWIDTH'b1111101100010100,
        `W_DATA_BITWIDTH'b0000000010010101,
        `W_DATA_BITWIDTH'b1111101001100110,
        `W_DATA_BITWIDTH'b1111101001100110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_DATA_BITWIDTH'b0000001011111110,
        `W_DATA_BITWIDTH'b0000000001111100,
        `W_DATA_BITWIDTH'b0000000100001101,
        `W_DATA_BITWIDTH'b0000001001111011,
        `W_DATA_BITWIDTH'b1111111011100110,
        `W_DATA_BITWIDTH'b1111111010000111,
        `W_DATA_BITWIDTH'b1111101111000001,
        `W_DATA_BITWIDTH'b1111111101100001,
        `W_DATA_BITWIDTH'b0000011011100110,
        `W_DATA_BITWIDTH'b0000000011100101,
        `W_DATA_BITWIDTH'b1111110011101111,
        `W_DATA_BITWIDTH'b0000000011101000,
        `W_DATA_BITWIDTH'b1111110100010101,
        `W_DATA_BITWIDTH'b1111110010010100,
        `W_DATA_BITWIDTH'b1111110011100001,
        `W_DATA_BITWIDTH'b0000000101010100,
        `W_DATA_BITWIDTH'b1111110111011100,
        `W_DATA_BITWIDTH'b1111110111011000,
        `W_DATA_BITWIDTH'b0000000101001100,
        `W_DATA_BITWIDTH'b1111110100010011,
        `W_DATA_BITWIDTH'b1111111010011111,
        `W_DATA_BITWIDTH'b0000001001100101,
        `W_DATA_BITWIDTH'b0000000111010101,
        `W_DATA_BITWIDTH'b1111100101110011,
        `W_DATA_BITWIDTH'b0000011010010111,
        `W_DATA_BITWIDTH'b0000000011000011,
        `W_DATA_BITWIDTH'b1111110101101010,
        `W_DATA_BITWIDTH'b0000000110111011,
        `W_DATA_BITWIDTH'b1111101110111011,
        `W_DATA_BITWIDTH'b0000010111100100,
        `W_DATA_BITWIDTH'b0000000110001111,
        `W_DATA_BITWIDTH'b0000010000001011,
        `W_DATA_BITWIDTH'b1111110111001100,
        `W_DATA_BITWIDTH'b1111111001100010,
        `W_DATA_BITWIDTH'b0000000101110101,
        `W_DATA_BITWIDTH'b1111101101101110,
        `W_DATA_BITWIDTH'b0000000100001110,
        `W_DATA_BITWIDTH'b0000000110111001,
        `W_DATA_BITWIDTH'b1111111100110110,
        `W_DATA_BITWIDTH'b1111111100101010,
        `W_DATA_BITWIDTH'b0000000111111111,
        `W_DATA_BITWIDTH'b0000100101101101,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110000000101,
        `W_DATA_BITWIDTH'b1111110000011011,
        `W_DATA_BITWIDTH'b0000000010110101,
        `W_DATA_BITWIDTH'b0000011010110011,
        `W_DATA_BITWIDTH'b1111111001101110,
        `W_DATA_BITWIDTH'b0000000101011110,
        `W_DATA_BITWIDTH'b1111111011001011,
        `W_DATA_BITWIDTH'b0000001101111000,
        `W_DATA_BITWIDTH'b0000011010000001,
        `W_DATA_BITWIDTH'b1111100010110110,
        `W_DATA_BITWIDTH'b1111110111010110,
        `W_DATA_BITWIDTH'b0000011010111110,
        `W_DATA_BITWIDTH'b1111101110100010,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b0000001000000110,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111100010100101,
        `W_DATA_BITWIDTH'b1111111011100000,
        `W_DATA_BITWIDTH'b0000001110100010,
        `W_DATA_BITWIDTH'b0000000111011111,
        `W_DATA_BITWIDTH'b1111110010111011,
        `W_DATA_BITWIDTH'b0000010000100101,
        `W_DATA_BITWIDTH'b0000010000100101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_DATA_BITWIDTH'b1111111101010101,
        `W_DATA_BITWIDTH'b0000000011101111,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110101011010,
        `W_DATA_BITWIDTH'b1111110101010100,
        `W_DATA_BITWIDTH'b0000001011110011,
        `W_DATA_BITWIDTH'b1111111001100101,
        `W_DATA_BITWIDTH'b0000010101111110,
        `W_DATA_BITWIDTH'b0000010010100101,
        `W_DATA_BITWIDTH'b1111011110010000,
        `W_DATA_BITWIDTH'b1111110001000001,
        `W_DATA_BITWIDTH'b0000001101001011,
        `W_DATA_BITWIDTH'b0000011001011010,
        `W_DATA_BITWIDTH'b1111100001111110,
        `W_DATA_BITWIDTH'b0000010010100111,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b1111111000111101,
        `W_DATA_BITWIDTH'b1111111011111100,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000110001000,
        `W_DATA_BITWIDTH'b1111110011001010,
        `W_DATA_BITWIDTH'b1111111001000011,
        `W_DATA_BITWIDTH'b1111111001011001,
        `W_DATA_BITWIDTH'b0000001010000101,
        `W_DATA_BITWIDTH'b0000001100001100,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111111001001011,
        `W_DATA_BITWIDTH'b0000010001001101,
        `W_DATA_BITWIDTH'b0000100000011111,
        `W_DATA_BITWIDTH'b1111100000100000,
        `W_DATA_BITWIDTH'b1111100111110111,
        `W_DATA_BITWIDTH'b0000001011100001,
        `W_DATA_BITWIDTH'b1111111101101011,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b0000001010100100,
        `W_DATA_BITWIDTH'b1111111000111110,
        `W_DATA_BITWIDTH'b0000001000000011,
        `W_DATA_BITWIDTH'b1111110101011011,
        `W_DATA_BITWIDTH'b1111111011010100,
        `W_DATA_BITWIDTH'b0000010010110001,
        `W_DATA_BITWIDTH'b1111110110001010,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b0000001110100101,
        `W_DATA_BITWIDTH'b0000000011100100,
        `W_DATA_BITWIDTH'b0000000111101001,
        `W_DATA_BITWIDTH'b0000001110011000,
        `W_DATA_BITWIDTH'b1111111101101010,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000001100101010,
        `W_DATA_BITWIDTH'b0000001001011111,
        `W_DATA_BITWIDTH'b1111111001010011,
        `W_DATA_BITWIDTH'b1111101010010111,
        `W_DATA_BITWIDTH'b1111110010010011,
        `W_DATA_BITWIDTH'b0000001111110100,
        `W_DATA_BITWIDTH'b0000000111011011,
        `W_DATA_BITWIDTH'b0000001011110101,
        `W_DATA_BITWIDTH'b1111100111101101,
        `W_DATA_BITWIDTH'b0000100000011000,
        `W_DATA_BITWIDTH'b1111111011111101,
        `W_DATA_BITWIDTH'b1111111011111101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_DATA_BITWIDTH'b1111110101111111,
        `W_DATA_BITWIDTH'b1111110101000101,
        `W_DATA_BITWIDTH'b0000001110111001,
        `W_DATA_BITWIDTH'b0000001100010101,
        `W_DATA_BITWIDTH'b1111110001010101,
        `W_DATA_BITWIDTH'b1111110110000011,
        `W_DATA_BITWIDTH'b1111110000110011,
        `W_DATA_BITWIDTH'b1111110011010001,
        `W_DATA_BITWIDTH'b0000001110101010,
        `W_DATA_BITWIDTH'b0000010000011111,
        `W_DATA_BITWIDTH'b1111110100011101,
        `W_DATA_BITWIDTH'b0000001010011111,
        `W_DATA_BITWIDTH'b0000001011001111,
        `W_DATA_BITWIDTH'b1111110110100001,
        `W_DATA_BITWIDTH'b1111101011111100,
        `W_DATA_BITWIDTH'b1111110110101110,
        `W_DATA_BITWIDTH'b0000001110000011,
        `W_DATA_BITWIDTH'b1111110000011010,
        `W_DATA_BITWIDTH'b0000001101101101,
        `W_DATA_BITWIDTH'b1111110101111010,
        `W_DATA_BITWIDTH'b1111110010101100,
        `W_DATA_BITWIDTH'b0000001011111000,
        `W_DATA_BITWIDTH'b1111110011100100,
        `W_DATA_BITWIDTH'b1111110100001011,
        `W_DATA_BITWIDTH'b1111110110001100,
        `W_DATA_BITWIDTH'b1111100111101010,
        `W_DATA_BITWIDTH'b1111110101001111,
        `W_DATA_BITWIDTH'b1111110011011100,
        `W_DATA_BITWIDTH'b1111110011010001,
        `W_DATA_BITWIDTH'b1111110111000100,
        `W_DATA_BITWIDTH'b0000001100001101,
        `W_DATA_BITWIDTH'b1111110111000100,
        `W_DATA_BITWIDTH'b0000001100010111,
        `W_DATA_BITWIDTH'b1111110000101111,
        `W_DATA_BITWIDTH'b1111100110110000,
        `W_DATA_BITWIDTH'b0000010111000111,
        `W_DATA_BITWIDTH'b0000001100100010,
        `W_DATA_BITWIDTH'b1111110001100110,
        `W_DATA_BITWIDTH'b1111110011000011,
        `W_DATA_BITWIDTH'b1111101111011111,
        `W_DATA_BITWIDTH'b1111101000111111,
        `W_DATA_BITWIDTH'b0000001011010011,
        `W_DATA_BITWIDTH'b0000001010011001,
        `W_DATA_BITWIDTH'b1111110011100111,
        `W_DATA_BITWIDTH'b0000001011011111,
        `W_DATA_BITWIDTH'b1111110110000101,
        `W_DATA_BITWIDTH'b0000010100001001,
        `W_DATA_BITWIDTH'b1111110110100100,
        `W_DATA_BITWIDTH'b0000010000011101,
        `W_DATA_BITWIDTH'b0000001010111011,
        `W_DATA_BITWIDTH'b1111100111110100,
        `W_DATA_BITWIDTH'b1111101010010100,
        `W_DATA_BITWIDTH'b0000010001010101,
        `W_DATA_BITWIDTH'b1111110110100100,
        `W_DATA_BITWIDTH'b1111101000100111,
        `W_DATA_BITWIDTH'b0000010100010001,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b0000001100110110,
        `W_DATA_BITWIDTH'b0000010010110000,
        `W_DATA_BITWIDTH'b1111110001100110,
        `W_DATA_BITWIDTH'b0000001100101000,
        `W_DATA_BITWIDTH'b1111110001011011,
        `W_DATA_BITWIDTH'b0000001011010001,
        `W_DATA_BITWIDTH'b0000011000001010,
        `W_DATA_BITWIDTH'b1111110011001011,
        `W_DATA_BITWIDTH'b1111110100111000,
        `W_DATA_BITWIDTH'b1111110011101100,
        `W_DATA_BITWIDTH'b1111110110110100,
        `W_DATA_BITWIDTH'b0000001100001000,
        `W_DATA_BITWIDTH'b0000001101111010,
        `W_DATA_BITWIDTH'b0000001100011100,
        `W_DATA_BITWIDTH'b1111110100000011,
        `W_DATA_BITWIDTH'b1111110101111100,
        `W_DATA_BITWIDTH'b1111101111101010,
        `W_DATA_BITWIDTH'b1111101100111011,
        `W_DATA_BITWIDTH'b1111110011100110,
        `W_DATA_BITWIDTH'b1111101010110101,
        `W_DATA_BITWIDTH'b1111101010110101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_DATA_BITWIDTH'b0000001101011111,
        `W_DATA_BITWIDTH'b0000010111001011,
        `W_DATA_BITWIDTH'b0000001111100110,
        `W_DATA_BITWIDTH'b0000010000111011,
        `W_DATA_BITWIDTH'b0000001110001001,
        `W_DATA_BITWIDTH'b1111101110111101,
        `W_DATA_BITWIDTH'b1111101010110101,
        `W_DATA_BITWIDTH'b1111101110000011,
        `W_DATA_BITWIDTH'b1111110110000011,
        `W_DATA_BITWIDTH'b1111110100110101,
        `W_DATA_BITWIDTH'b1111110101011001,
        `W_DATA_BITWIDTH'b0000001111001011,
        `W_DATA_BITWIDTH'b1111110110100111,
        `W_DATA_BITWIDTH'b1111110100101010,
        `W_DATA_BITWIDTH'b1111110010100000,
        `W_DATA_BITWIDTH'b1111101111100000,
        `W_DATA_BITWIDTH'b0000010010100100,
        `W_DATA_BITWIDTH'b0000001101101100,
        `W_DATA_BITWIDTH'b0000001001011011,
        `W_DATA_BITWIDTH'b1111110101011110,
        `W_DATA_BITWIDTH'b1111110010110001,
        `W_DATA_BITWIDTH'b1111101111101101,
        `W_DATA_BITWIDTH'b0000001100100001,
        `W_DATA_BITWIDTH'b0000001111001011,
        `W_DATA_BITWIDTH'b0000001011000110,
        `W_DATA_BITWIDTH'b1111101101011101,
        `W_DATA_BITWIDTH'b0000001010010011,
        `W_DATA_BITWIDTH'b1111110000000000,
        `W_DATA_BITWIDTH'b0000001001111100,
        `W_DATA_BITWIDTH'b0000001011010101,
        `W_DATA_BITWIDTH'b1111110011111011,
        `W_DATA_BITWIDTH'b1111101110011001,
        `W_DATA_BITWIDTH'b1111110110001000,
        `W_DATA_BITWIDTH'b0000001000111101,
        `W_DATA_BITWIDTH'b1111110110111111,
        `W_DATA_BITWIDTH'b0000001001011001,
        `W_DATA_BITWIDTH'b0000001010101100,
        `W_DATA_BITWIDTH'b1111110010110101,
        `W_DATA_BITWIDTH'b0000001000111100,
        `W_DATA_BITWIDTH'b1111110100100010,
        `W_DATA_BITWIDTH'b1111110001110100,
        `W_DATA_BITWIDTH'b1111101101011011,
        `W_DATA_BITWIDTH'b1111110101100010,
        `W_DATA_BITWIDTH'b1111110101101110,
        `W_DATA_BITWIDTH'b1111110101100101,
        `W_DATA_BITWIDTH'b0000001001111101,
        `W_DATA_BITWIDTH'b1111110100001100,
        `W_DATA_BITWIDTH'b0000010000011100,
        `W_DATA_BITWIDTH'b1111110101111001,
        `W_DATA_BITWIDTH'b0000001101100011,
        `W_DATA_BITWIDTH'b1111110101010010,
        `W_DATA_BITWIDTH'b1111110110101111,
        `W_DATA_BITWIDTH'b1111110101100110,
        `W_DATA_BITWIDTH'b1111110101100111,
        `W_DATA_BITWIDTH'b0000001100101110,
        `W_DATA_BITWIDTH'b0000001011100111,
        `W_DATA_BITWIDTH'b1111110010110011,
        `W_DATA_BITWIDTH'b0000010101110101,
        `W_DATA_BITWIDTH'b0000001001011111,
        `W_DATA_BITWIDTH'b1111100101101101,
        `W_DATA_BITWIDTH'b1111110100010010,
        `W_DATA_BITWIDTH'b0000001110100000,
        `W_DATA_BITWIDTH'b1111110011101110,
        `W_DATA_BITWIDTH'b1111110010110100,
        `W_DATA_BITWIDTH'b1111101111110101,
        `W_DATA_BITWIDTH'b1111101010010001,
        `W_DATA_BITWIDTH'b0000010010001110,
        `W_DATA_BITWIDTH'b0000001101011111,
        `W_DATA_BITWIDTH'b1111101000100110,
        `W_DATA_BITWIDTH'b1111110101010111,
        `W_DATA_BITWIDTH'b0000001001010010,
        `W_DATA_BITWIDTH'b0000001001111010,
        `W_DATA_BITWIDTH'b1111110101110001,
        `W_DATA_BITWIDTH'b0000001111011011,
        `W_DATA_BITWIDTH'b0000001111011011,
        `W_DATA_BITWIDTH'b0000001101101001,
        `W_DATA_BITWIDTH'b0000010010001000,
        `W_DATA_BITWIDTH'b0000001010011001,
        `W_DATA_BITWIDTH'b0000001011000011,
        `W_DATA_BITWIDTH'b0000001100001010,
        `W_DATA_BITWIDTH'b1111110100110010,
        `W_DATA_BITWIDTH'b1111110100110100,
        `W_DATA_BITWIDTH'b1111110100101100,
        `W_DATA_BITWIDTH'b1111110100100111,
        `W_DATA_BITWIDTH'b0000001100010010,
        `W_DATA_BITWIDTH'b0000001100010010
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_DATA_BITWIDTH'b1111110101111000,
        `W_DATA_BITWIDTH'b0000001100011110,
        `W_DATA_BITWIDTH'b0000001111111111,
        `W_DATA_BITWIDTH'b1111110011111001,
        `W_DATA_BITWIDTH'b1111110110000100,
        `W_DATA_BITWIDTH'b1111101111000110,
        `W_DATA_BITWIDTH'b1111110110010110,
        `W_DATA_BITWIDTH'b1111110000101110,
        `W_DATA_BITWIDTH'b0000010001010110,
        `W_DATA_BITWIDTH'b1111101010001110,
        `W_DATA_BITWIDTH'b0000010000001111,
        `W_DATA_BITWIDTH'b1111101111100111,
        `W_DATA_BITWIDTH'b0000001000111011,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b1111110101011011,
        `W_DATA_BITWIDTH'b1111110011100001,
        `W_DATA_BITWIDTH'b1111110011010111,
        `W_DATA_BITWIDTH'b1111110001101011,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b1111110000101010,
        `W_DATA_BITWIDTH'b1111110101010010,
        `W_DATA_BITWIDTH'b0000010001000110,
        `W_DATA_BITWIDTH'b1111101111001110,
        `W_DATA_BITWIDTH'b0000001011110001,
        `W_DATA_BITWIDTH'b0000001100011001,
        `W_DATA_BITWIDTH'b1111110011000110,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b0000010000000100,
        `W_DATA_BITWIDTH'b1111110101001100,
        `W_DATA_BITWIDTH'b1111110111000010,
        `W_DATA_BITWIDTH'b0000001110110101,
        `W_DATA_BITWIDTH'b1111101110001100,
        `W_DATA_BITWIDTH'b1111110010000111,
        `W_DATA_BITWIDTH'b0000001010111010,
        `W_DATA_BITWIDTH'b1111110100110110,
        `W_DATA_BITWIDTH'b1111110000110010,
        `W_DATA_BITWIDTH'b1111110011101110,
        `W_DATA_BITWIDTH'b1111101101101000,
        `W_DATA_BITWIDTH'b1111110011110101,
        `W_DATA_BITWIDTH'b0000010100111111,
        `W_DATA_BITWIDTH'b1111101111101011,
        `W_DATA_BITWIDTH'b1111110001001100,
        `W_DATA_BITWIDTH'b0000011010110011,
        `W_DATA_BITWIDTH'b0000010011111011,
        `W_DATA_BITWIDTH'b0000001100010001,
        `W_DATA_BITWIDTH'b0000011011000000,
        `W_DATA_BITWIDTH'b1111101001110000,
        `W_DATA_BITWIDTH'b1111110110011111,
        `W_DATA_BITWIDTH'b1111110000101010,
        `W_DATA_BITWIDTH'b1111110011110011,
        `W_DATA_BITWIDTH'b0000001010111101,
        `W_DATA_BITWIDTH'b1111100100101101,
        `W_DATA_BITWIDTH'b1111110100001110,
        `W_DATA_BITWIDTH'b1111110110111111,
        `W_DATA_BITWIDTH'b1111101000010110,
        `W_DATA_BITWIDTH'b0000010001011111,
        `W_DATA_BITWIDTH'b1111110010101101,
        `W_DATA_BITWIDTH'b0000010010101011,
        `W_DATA_BITWIDTH'b0000001001100111,
        `W_DATA_BITWIDTH'b1111101011111101,
        `W_DATA_BITWIDTH'b1111110110100010,
        `W_DATA_BITWIDTH'b0000001001000101,
        `W_DATA_BITWIDTH'b1111110100101101,
        `W_DATA_BITWIDTH'b0000001001001011,
        `W_DATA_BITWIDTH'b1111110010001011,
        `W_DATA_BITWIDTH'b1111110010001011
    };

// w_data
