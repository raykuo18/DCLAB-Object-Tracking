`include "header.h"

module Top(
	input              i_clk,
	input              i_rst_n,
	input              i_start,
	output logic [3:0] o_random_out
);
    // ========================== Parameters definition ==================================

        // ----- WMem --------
            // w_data
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
                '{
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b1111110111110001,
                    `W_DATA_BITWIDTH'b0000000010111001,
                    `W_DATA_BITWIDTH'b1111111001001000,
                    `W_DATA_BITWIDTH'b1111111100101100,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000001011101001,
                    `W_DATA_BITWIDTH'b0000001110000101,
                    `W_DATA_BITWIDTH'b1111100101001100,
                    `W_DATA_BITWIDTH'b1111101000011010,
                    `W_DATA_BITWIDTH'b0000001000111111,
                    `W_DATA_BITWIDTH'b1111011110101000,
                    `W_DATA_BITWIDTH'b1111111011101100,
                    `W_DATA_BITWIDTH'b0000110100100001,
                    `W_DATA_BITWIDTH'b0000011110000000,
                    `W_DATA_BITWIDTH'b1111011101111100,
                    `W_DATA_BITWIDTH'b0000101111111011,
                    `W_DATA_BITWIDTH'b1111110110101010,
                    `W_DATA_BITWIDTH'b0000010000001010,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b1111001101110010,
                    `W_DATA_BITWIDTH'b0000101101101000,
                    `W_DATA_BITWIDTH'b0000001101100100,
                    `W_DATA_BITWIDTH'b0000100001011110,
                    `W_DATA_BITWIDTH'b1111101101101010,
                    `W_DATA_BITWIDTH'b0000010110010101,
                    `W_DATA_BITWIDTH'b0000100011000111,
                    `W_DATA_BITWIDTH'b1111111001000000,
                    `W_DATA_BITWIDTH'b1111101000010001,
                    `W_DATA_BITWIDTH'b0000000111110100,
                    `W_DATA_BITWIDTH'b0000001111001101,
                    `W_DATA_BITWIDTH'b0000100001011110,
                    `W_DATA_BITWIDTH'b0000010110100100,
                    `W_DATA_BITWIDTH'b0000001001101110,
                    `W_DATA_BITWIDTH'b1111110000000001,
                    `W_DATA_BITWIDTH'b1111100111111011,
                    `W_DATA_BITWIDTH'b1111101010101100,
                    `W_DATA_BITWIDTH'b1111011110100100,
                    `W_DATA_BITWIDTH'b0000011011011001,
                    `W_DATA_BITWIDTH'b1111101111111110,
                    `W_DATA_BITWIDTH'b0000010000110000,
                    `W_DATA_BITWIDTH'b1111110110111010,
                    `W_DATA_BITWIDTH'b1111100011101101,
                    `W_DATA_BITWIDTH'b1111110010001101,
                    `W_DATA_BITWIDTH'b0000001110100011,
                    `W_DATA_BITWIDTH'b0000011111010101,
                    `W_DATA_BITWIDTH'b1111101110111101,
                    `W_DATA_BITWIDTH'b0000010101111100,
                    `W_DATA_BITWIDTH'b0000001011110110,
                    `W_DATA_BITWIDTH'b0000010010100011,
                    `W_DATA_BITWIDTH'b0000000100100010,
                    `W_DATA_BITWIDTH'b0000010110111000,
                    `W_DATA_BITWIDTH'b0000000100101001,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000111000001,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111001101111,
                    `W_DATA_BITWIDTH'b1111111000010110,
                    `W_DATA_BITWIDTH'b0000000111101010,
                    `W_DATA_BITWIDTH'b0000000111001111,
                    `W_DATA_BITWIDTH'b1111110101100100,
                    `W_DATA_BITWIDTH'b0000010001001100,
                    `W_DATA_BITWIDTH'b0000010010000011,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000100101011,
                    `W_DATA_BITWIDTH'b0000001001100011,
                    `W_DATA_BITWIDTH'b1111101111010111,
                    `W_DATA_BITWIDTH'b1111101010110111,
                    `W_DATA_BITWIDTH'b0000001111100111,
                    `W_DATA_BITWIDTH'b0000001101000010,
                    `W_DATA_BITWIDTH'b1111101110111001,
                    `W_DATA_BITWIDTH'b0000010010101110,
                    `W_DATA_BITWIDTH'b0000001111100110,
                    `W_DATA_BITWIDTH'b0000010010010110,
                    `W_DATA_BITWIDTH'b1111110100101101,
                    `W_DATA_BITWIDTH'b1111111011010101,
                    `W_DATA_BITWIDTH'b1111110100001000,
                    `W_DATA_BITWIDTH'b1111111011001011,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111010100111,
                    `W_DATA_BITWIDTH'b1111111001011111,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111110101010000,
                    `W_DATA_BITWIDTH'b1111111001001110,
                    `W_DATA_BITWIDTH'b1111101010011110,
                    `W_DATA_BITWIDTH'b1111100100101111,
                    `W_DATA_BITWIDTH'b1111110010101000,
                    `W_DATA_BITWIDTH'b1111010110111011,
                    `W_DATA_BITWIDTH'b0000001011110000,
                    `W_DATA_BITWIDTH'b1111110010011011,
                    `W_DATA_BITWIDTH'b0000000111101001,
                    `W_DATA_BITWIDTH'b0000001101010010,
                    `W_DATA_BITWIDTH'b0000000010011101,
                    `W_DATA_BITWIDTH'b1111111000010111,
                    `W_DATA_BITWIDTH'b0000011110111111,
                    `W_DATA_BITWIDTH'b0000100010111000,
                    `W_DATA_BITWIDTH'b0000001000011010,
                    `W_DATA_BITWIDTH'b1111100110001010,
                    `W_DATA_BITWIDTH'b1111110011110100,
                    `W_DATA_BITWIDTH'b1111101011111011,
                    `W_DATA_BITWIDTH'b0000001011001011,
                    `W_DATA_BITWIDTH'b0000001000110010,
                    `W_DATA_BITWIDTH'b1111110010001011,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b1111111101111110,
                    `W_DATA_BITWIDTH'b0000001001111101,
                    `W_DATA_BITWIDTH'b0000001000001111,
                    `W_DATA_BITWIDTH'b1111110111000001,
                    `W_DATA_BITWIDTH'b1111101000000010,
                    `W_DATA_BITWIDTH'b0000010000001111,
                    `W_DATA_BITWIDTH'b1111110101010001,
                    `W_DATA_BITWIDTH'b0000000101110110,
                    `W_DATA_BITWIDTH'b0000001100010100,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b0000000110000101,
                    `W_DATA_BITWIDTH'b1111111100111100,
                    `W_DATA_BITWIDTH'b0000001000011100,
                    `W_DATA_BITWIDTH'b0000001000110011,
                    `W_DATA_BITWIDTH'b0000000110011001,
                    `W_DATA_BITWIDTH'b0000000101111100,
                    `W_DATA_BITWIDTH'b0000001001100000,
                    `W_DATA_BITWIDTH'b1111110110110110,
                    `W_DATA_BITWIDTH'b1111110110110110
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000101011111,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b0000000111100111,
                    `W_DATA_BITWIDTH'b0000000100101110,
                    `W_DATA_BITWIDTH'b0000001000110010,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b1111110111110110,
                    `W_DATA_BITWIDTH'b1111100111000001,
                    `W_DATA_BITWIDTH'b1111110111010101,
                    `W_DATA_BITWIDTH'b1111110000111010,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b0000000011011000,
                    `W_DATA_BITWIDTH'b1111111010010100,
                    `W_DATA_BITWIDTH'b0000000101001111,
                    `W_DATA_BITWIDTH'b1111101100011101,
                    `W_DATA_BITWIDTH'b0000010110011010,
                    `W_DATA_BITWIDTH'b1111110100111010,
                    `W_DATA_BITWIDTH'b1111100010111110,
                    `W_DATA_BITWIDTH'b1111011101011101,
                    `W_DATA_BITWIDTH'b1111011000001011,
                    `W_DATA_BITWIDTH'b1111110101001011,
                    `W_DATA_BITWIDTH'b0000010111101111,
                    `W_DATA_BITWIDTH'b1111111000000100,
                    `W_DATA_BITWIDTH'b0000101110010000,
                    `W_DATA_BITWIDTH'b1111011100111010,
                    `W_DATA_BITWIDTH'b0000001101111000,
                    `W_DATA_BITWIDTH'b1111101010101101,
                    `W_DATA_BITWIDTH'b0000100000101000,
                    `W_DATA_BITWIDTH'b0000101110110101,
                    `W_DATA_BITWIDTH'b1111101100111000,
                    `W_DATA_BITWIDTH'b1111101100011100,
                    `W_DATA_BITWIDTH'b1111011100100010,
                    `W_DATA_BITWIDTH'b0000100000110000,
                    `W_DATA_BITWIDTH'b0000011110000000,
                    `W_DATA_BITWIDTH'b0000011000010101,
                    `W_DATA_BITWIDTH'b0000001010000011,
                    `W_DATA_BITWIDTH'b0000010000010000,
                    `W_DATA_BITWIDTH'b0000000011111110,
                    `W_DATA_BITWIDTH'b1111101100111110,
                    `W_DATA_BITWIDTH'b1111101110110110,
                    `W_DATA_BITWIDTH'b0000001000100110,
                    `W_DATA_BITWIDTH'b0000010011101111,
                    `W_DATA_BITWIDTH'b0000001010110001,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b1111100011110100,
                    `W_DATA_BITWIDTH'b1111100110101001,
                    `W_DATA_BITWIDTH'b0000011101011110,
                    `W_DATA_BITWIDTH'b1111111011101000,
                    `W_DATA_BITWIDTH'b0000001110110001,
                    `W_DATA_BITWIDTH'b0000001101001111,
                    `W_DATA_BITWIDTH'b0000001110100111,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b1111101000011110,
                    `W_DATA_BITWIDTH'b1111100110000110,
                    `W_DATA_BITWIDTH'b0000000111110100,
                    `W_DATA_BITWIDTH'b1111101011101001,
                    `W_DATA_BITWIDTH'b1111111011010000,
                    `W_DATA_BITWIDTH'b0000011100111011,
                    `W_DATA_BITWIDTH'b1111111001010001,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000100001001,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b1111111010010000,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000110101011,
                    `W_DATA_BITWIDTH'b0000000011001110,
                    `W_DATA_BITWIDTH'b0000001011100010,
                    `W_DATA_BITWIDTH'b1111111001100000,
                    `W_DATA_BITWIDTH'b0000010000010010,
                    `W_DATA_BITWIDTH'b0000000100000100,
                    `W_DATA_BITWIDTH'b1111111011101001,
                    `W_DATA_BITWIDTH'b1111101101101001,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111111100100110,
                    `W_DATA_BITWIDTH'b1111110011011001,
                    `W_DATA_BITWIDTH'b1111110011110101,
                    `W_DATA_BITWIDTH'b0000000110111011,
                    `W_DATA_BITWIDTH'b0000001000110011,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b0000010010110111,
                    `W_DATA_BITWIDTH'b0000001000010010,
                    `W_DATA_BITWIDTH'b0000001111100010,
                    `W_DATA_BITWIDTH'b1111101110000101,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b0000000100011110,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b1111101111111100,
                    `W_DATA_BITWIDTH'b0000100011111111,
                    `W_DATA_BITWIDTH'b0000001001011111,
                    `W_DATA_BITWIDTH'b1111011100110011,
                    `W_DATA_BITWIDTH'b0000000101111010,
                    `W_DATA_BITWIDTH'b0000100001010011,
                    `W_DATA_BITWIDTH'b0000100100011011,
                    `W_DATA_BITWIDTH'b1111100011111100,
                    `W_DATA_BITWIDTH'b0000000011100010,
                    `W_DATA_BITWIDTH'b0000000110001010,
                    `W_DATA_BITWIDTH'b0000000101101101,
                    `W_DATA_BITWIDTH'b0000000100110111,
                    `W_DATA_BITWIDTH'b1111110000110011,
                    `W_DATA_BITWIDTH'b1111110011001100,
                    `W_DATA_BITWIDTH'b0000010011110100,
                    `W_DATA_BITWIDTH'b1111100001111001,
                    `W_DATA_BITWIDTH'b1111101011000000,
                    `W_DATA_BITWIDTH'b0000011000110100,
                    `W_DATA_BITWIDTH'b1111111000010010,
                    `W_DATA_BITWIDTH'b1111110101110110,
                    `W_DATA_BITWIDTH'b1111110000001110,
                    `W_DATA_BITWIDTH'b1111110101100100,
                    `W_DATA_BITWIDTH'b0000001110111111,
                    `W_DATA_BITWIDTH'b1111111101110011,
                    `W_DATA_BITWIDTH'b0000000111101110,
                    `W_DATA_BITWIDTH'b0000001100100011,
                    `W_DATA_BITWIDTH'b1111110110110100,
                    `W_DATA_BITWIDTH'b1111111100110101,
                    `W_DATA_BITWIDTH'b0000000111111110,
                    `W_DATA_BITWIDTH'b0000001101111010,
                    `W_DATA_BITWIDTH'b1111111000111010,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b1111110010000001,
                    `W_DATA_BITWIDTH'b1111110000111011,
                    `W_DATA_BITWIDTH'b1111110110111010,
                    `W_DATA_BITWIDTH'b1111111001000010,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b1111110111110111,
                    `W_DATA_BITWIDTH'b0000000111000111,
                    `W_DATA_BITWIDTH'b0000001011100000,
                    `W_DATA_BITWIDTH'b0000000101101011,
                    `W_DATA_BITWIDTH'b0000000101101011
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b1111111001101101,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000101101111,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b0000000110001110,
                    `W_DATA_BITWIDTH'b0000000111000011,
                    `W_DATA_BITWIDTH'b0000000100111000,
                    `W_DATA_BITWIDTH'b0000001010100011,
                    `W_DATA_BITWIDTH'b0000011001010111,
                    `W_DATA_BITWIDTH'b0000010111100000,
                    `W_DATA_BITWIDTH'b1111110101010110,
                    `W_DATA_BITWIDTH'b0000001110110110,
                    `W_DATA_BITWIDTH'b0000010000001100,
                    `W_DATA_BITWIDTH'b0000011101011110,
                    `W_DATA_BITWIDTH'b0000100011000010,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b0000010110101000,
                    `W_DATA_BITWIDTH'b1111110111000001,
                    `W_DATA_BITWIDTH'b1111101101110010,
                    `W_DATA_BITWIDTH'b1111100001100100,
                    `W_DATA_BITWIDTH'b1111011100010000,
                    `W_DATA_BITWIDTH'b0000001010010010,
                    `W_DATA_BITWIDTH'b0000100010011111,
                    `W_DATA_BITWIDTH'b1111111001101100,
                    `W_DATA_BITWIDTH'b1111100000100001,
                    `W_DATA_BITWIDTH'b1111110001100011,
                    `W_DATA_BITWIDTH'b1111110101110110,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b1111011101000001,
                    `W_DATA_BITWIDTH'b1111011110011101,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b0000001110110100,
                    `W_DATA_BITWIDTH'b1111101101011100,
                    `W_DATA_BITWIDTH'b0000000110010011,
                    `W_DATA_BITWIDTH'b1111101000101111,
                    `W_DATA_BITWIDTH'b1111111001100001,
                    `W_DATA_BITWIDTH'b1111110000101001,
                    `W_DATA_BITWIDTH'b1111101101110000,
                    `W_DATA_BITWIDTH'b0000001101010011,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000010011110101,
                    `W_DATA_BITWIDTH'b1111100010100000,
                    `W_DATA_BITWIDTH'b1111011000000110,
                    `W_DATA_BITWIDTH'b1111101001101111,
                    `W_DATA_BITWIDTH'b1111110101000000,
                    `W_DATA_BITWIDTH'b0000001011000000,
                    `W_DATA_BITWIDTH'b0000011010001000,
                    `W_DATA_BITWIDTH'b0000001000110001,
                    `W_DATA_BITWIDTH'b0000010111001000,
                    `W_DATA_BITWIDTH'b1111101010011000,
                    `W_DATA_BITWIDTH'b1111100001101011,
                    `W_DATA_BITWIDTH'b1111111011001100,
                    `W_DATA_BITWIDTH'b1111100010111100,
                    `W_DATA_BITWIDTH'b0000001110101000,
                    `W_DATA_BITWIDTH'b0000000100011011,
                    `W_DATA_BITWIDTH'b0000011111001100,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b0000000101100011,
                    `W_DATA_BITWIDTH'b1111111011001101,
                    `W_DATA_BITWIDTH'b0000001001000110,
                    `W_DATA_BITWIDTH'b0000001001000011,
                    `W_DATA_BITWIDTH'b1111111011101110,
                    `W_DATA_BITWIDTH'b0000001110000101,
                    `W_DATA_BITWIDTH'b0000001110011101,
                    `W_DATA_BITWIDTH'b1111111000001111,
                    `W_DATA_BITWIDTH'b0000001011110001,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b0000000100100001,
                    `W_DATA_BITWIDTH'b0000001011111111,
                    `W_DATA_BITWIDTH'b1111110101010110,
                    `W_DATA_BITWIDTH'b1111111011100001,
                    `W_DATA_BITWIDTH'b1111101101010001,
                    `W_DATA_BITWIDTH'b1111110001110111,
                    `W_DATA_BITWIDTH'b0000001010111101,
                    `W_DATA_BITWIDTH'b1111110001101001,
                    `W_DATA_BITWIDTH'b0000001010100110,
                    `W_DATA_BITWIDTH'b0000001101010001,
                    `W_DATA_BITWIDTH'b1111110001001111,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b1111111011100110,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b0000000101000111,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b0000010111010101,
                    `W_DATA_BITWIDTH'b0000011011111100,
                    `W_DATA_BITWIDTH'b0000011010010110,
                    `W_DATA_BITWIDTH'b0000001000100010,
                    `W_DATA_BITWIDTH'b1111101010000010,
                    `W_DATA_BITWIDTH'b1111111000101001,
                    `W_DATA_BITWIDTH'b1111110110010100,
                    `W_DATA_BITWIDTH'b0000000111011110,
                    `W_DATA_BITWIDTH'b1111101011011110,
                    `W_DATA_BITWIDTH'b0000011111111101,
                    `W_DATA_BITWIDTH'b1111011101110110,
                    `W_DATA_BITWIDTH'b1111110111011101,
                    `W_DATA_BITWIDTH'b1111111000101110,
                    `W_DATA_BITWIDTH'b0000010011001111,
                    `W_DATA_BITWIDTH'b0000001010011000,
                    `W_DATA_BITWIDTH'b1111101011100110,
                    `W_DATA_BITWIDTH'b1111111000011100,
                    `W_DATA_BITWIDTH'b1111111000010110,
                    `W_DATA_BITWIDTH'b1111110101011010,
                    `W_DATA_BITWIDTH'b1111110101001001,
                    `W_DATA_BITWIDTH'b1111111001100010,
                    `W_DATA_BITWIDTH'b0000000110110101,
                    `W_DATA_BITWIDTH'b0000000110111010,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b0000001011100010,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b0000001010000000,
                    `W_DATA_BITWIDTH'b1111111001011011,
                    `W_DATA_BITWIDTH'b1111111011011111,
                    `W_DATA_BITWIDTH'b1111110001101000,
                    `W_DATA_BITWIDTH'b1111110111010101,
                    `W_DATA_BITWIDTH'b1111111010100010,
                    `W_DATA_BITWIDTH'b1111111001011001,
                    `W_DATA_BITWIDTH'b1111111001111110,
                    `W_DATA_BITWIDTH'b0000001010101001,
                    `W_DATA_BITWIDTH'b1111111001011110,
                    `W_DATA_BITWIDTH'b0000000100010001,
                    `W_DATA_BITWIDTH'b1111111000010110,
                    `W_DATA_BITWIDTH'b1111111000010110
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111111101101010,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111001010010,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b0000000010011101,
                    `W_DATA_BITWIDTH'b1111111011010101,
                    `W_DATA_BITWIDTH'b0000000011011001,
                    `W_DATA_BITWIDTH'b0000000100110100,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000010010010,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b0000000110001101,
                    `W_DATA_BITWIDTH'b1111111010111110,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b1111111101001111,
                    `W_DATA_BITWIDTH'b0000000101001001,
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b0000000010001000,
                    `W_DATA_BITWIDTH'b1111111101001110,
                    `W_DATA_BITWIDTH'b1111111100000100,
                    `W_DATA_BITWIDTH'b0000000010111100,
                    `W_DATA_BITWIDTH'b0000000011101000,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b1111111011100111,
                    `W_DATA_BITWIDTH'b1111111101101001,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111100001000,
                    `W_DATA_BITWIDTH'b0000000011000010,
                    `W_DATA_BITWIDTH'b0000000010100100,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b1111111011000111,
                    `W_DATA_BITWIDTH'b0000000011000000,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b1111111001110100,
                    `W_DATA_BITWIDTH'b1111111001000101,
                    `W_DATA_BITWIDTH'b0000000100111001,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b0000000110001111,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b0000000101100010,
                    `W_DATA_BITWIDTH'b1111111100001101,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111011010110,
                    `W_DATA_BITWIDTH'b0000000011011101,
                    `W_DATA_BITWIDTH'b1111110111000000,
                    `W_DATA_BITWIDTH'b1111111001011011,
                    `W_DATA_BITWIDTH'b1111111000101101,
                    `W_DATA_BITWIDTH'b0000000100101110,
                    `W_DATA_BITWIDTH'b0000000011100011,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111110111110011,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b1111111101011101,
                    `W_DATA_BITWIDTH'b0000000100010011,
                    `W_DATA_BITWIDTH'b1111111011011000,
                    `W_DATA_BITWIDTH'b1111111101000011,
                    `W_DATA_BITWIDTH'b1111111101000110,
                    `W_DATA_BITWIDTH'b0000000100010110,
                    `W_DATA_BITWIDTH'b0000000011100001,
                    `W_DATA_BITWIDTH'b1111111011011010,
                    `W_DATA_BITWIDTH'b1111110111011001,
                    `W_DATA_BITWIDTH'b1111111010110110,
                    `W_DATA_BITWIDTH'b1111111011001010,
                    `W_DATA_BITWIDTH'b0000000100001011,
                    `W_DATA_BITWIDTH'b0000000010010100,
                    `W_DATA_BITWIDTH'b1111111011001110,
                    `W_DATA_BITWIDTH'b1111111001100010,
                    `W_DATA_BITWIDTH'b0000000010100101,
                    `W_DATA_BITWIDTH'b1111111010101110,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b1111111010101000,
                    `W_DATA_BITWIDTH'b1111111100111001,
                    `W_DATA_BITWIDTH'b1111111010110010,
                    `W_DATA_BITWIDTH'b0000000010110101,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111100011100,
                    `W_DATA_BITWIDTH'b1111110110001010,
                    `W_DATA_BITWIDTH'b0000000010110111,
                    `W_DATA_BITWIDTH'b0000000111001000,
                    `W_DATA_BITWIDTH'b0000000100101101,
                    `W_DATA_BITWIDTH'b1111111010111001,
                    `W_DATA_BITWIDTH'b0000000011001101,
                    `W_DATA_BITWIDTH'b1111110001110111,
                    `W_DATA_BITWIDTH'b1111111000100001,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b1111110100001001,
                    `W_DATA_BITWIDTH'b1111111010010111,
                    `W_DATA_BITWIDTH'b1111110111001110,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b1111111001001100,
                    `W_DATA_BITWIDTH'b1111110110100001,
                    `W_DATA_BITWIDTH'b1111111011010010,
                    `W_DATA_BITWIDTH'b0000000101110000,
                    `W_DATA_BITWIDTH'b1111111010111010,
                    `W_DATA_BITWIDTH'b1111111011101010,
                    `W_DATA_BITWIDTH'b1111111010100011,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111100100101,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b1111111011011011,
                    `W_DATA_BITWIDTH'b0000000100110100,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b0000000011010111,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b1111111101100000,
                    `W_DATA_BITWIDTH'b0000000010110010,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b0000000100101110,
                    `W_DATA_BITWIDTH'b0000000010100000,
                    `W_DATA_BITWIDTH'b1111111010010101,
                    `W_DATA_BITWIDTH'b1111111101001100,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b1111111010110101,
                    `W_DATA_BITWIDTH'b1111111101111100,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b1111111100110111,
                    `W_DATA_BITWIDTH'b1111111011011100,
                    `W_DATA_BITWIDTH'b1111111100001011,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111100101110,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b1111111011110000,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b0000000100100101,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b1111111010100010,
                    `W_DATA_BITWIDTH'b1111111010110000,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b0000000011010000,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b0000000011000010,
                    `W_DATA_BITWIDTH'b0000000100001101,
                    `W_DATA_BITWIDTH'b0000000011101101,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b1111111011101101,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b1111111101011110,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b0000000101001001,
                    `W_DATA_BITWIDTH'b0000000011000000,
                    `W_DATA_BITWIDTH'b0000000101110110,
                    `W_DATA_BITWIDTH'b0000000010110110,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b0000000011010011,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111111100100010,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000011100001,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b1111111101001001,
                    `W_DATA_BITWIDTH'b1111111101010001,
                    `W_DATA_BITWIDTH'b1111111101100101,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111100001011,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000011100011,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b1111111010101110,
                    `W_DATA_BITWIDTH'b1111111011000011,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b1111111011010011,
                    `W_DATA_BITWIDTH'b1111111101000000,
                    `W_DATA_BITWIDTH'b1111111001111100,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b0000000011101000,
                    `W_DATA_BITWIDTH'b1111111101101111,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b0000000010111001,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000100010010,
                    `W_DATA_BITWIDTH'b0000000100110100,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b1111111010110110,
                    `W_DATA_BITWIDTH'b1111111100111110,
                    `W_DATA_BITWIDTH'b0000000100001010,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b0000000101111001,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111011101110,
                    `W_DATA_BITWIDTH'b0000000101111101,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111010100011,
                    `W_DATA_BITWIDTH'b0000000100100011,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b1111110110111010,
                    `W_DATA_BITWIDTH'b1111111101000110,
                    `W_DATA_BITWIDTH'b1111111011001000,
                    `W_DATA_BITWIDTH'b0000000011010001,
                    `W_DATA_BITWIDTH'b1111110001011000,
                    `W_DATA_BITWIDTH'b1111111100000100,
                    `W_DATA_BITWIDTH'b0000000111001101,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b0000000101001011,
                    `W_DATA_BITWIDTH'b0000000110110111,
                    `W_DATA_BITWIDTH'b1111110101001010,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000001000010101,
                    `W_DATA_BITWIDTH'b1111111001010010,
                    `W_DATA_BITWIDTH'b0000000110001000,
                    `W_DATA_BITWIDTH'b0000000011100110,
                    `W_DATA_BITWIDTH'b1111110111000110,
                    `W_DATA_BITWIDTH'b1111111001101001,
                    `W_DATA_BITWIDTH'b1111111001110011,
                    `W_DATA_BITWIDTH'b1111111101001010,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b0000000101010010,
                    `W_DATA_BITWIDTH'b0000000100101000,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b1111111001111100,
                    `W_DATA_BITWIDTH'b1111111100000011,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b0000000110001101,
                    `W_DATA_BITWIDTH'b1111111101001011,
                    `W_DATA_BITWIDTH'b1111111010111110,
                    `W_DATA_BITWIDTH'b1111111001100101,
                    `W_DATA_BITWIDTH'b0000001000110111,
                    `W_DATA_BITWIDTH'b1111111000100010,
                    `W_DATA_BITWIDTH'b1111111100011001,
                    `W_DATA_BITWIDTH'b0000001001000111,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b1111111101111100,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111100101010,
                    `W_DATA_BITWIDTH'b0000000010010100,
                    `W_DATA_BITWIDTH'b1111111100101010,
                    `W_DATA_BITWIDTH'b1111111101010010,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111111101011100,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b1111111100010100,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b1111111011001110,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000100001101,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b1111111101011100,
                    `W_DATA_BITWIDTH'b0000000101100010,
                    `W_DATA_BITWIDTH'b0000000011001001,
                    `W_DATA_BITWIDTH'b1111111011100101,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000011100010,
                    `W_DATA_BITWIDTH'b0000000100011100,
                    `W_DATA_BITWIDTH'b1111111011100111,
                    `W_DATA_BITWIDTH'b0000000110000011,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b1111111011110010,
                    `W_DATA_BITWIDTH'b1111111100101110,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b1111111000010001,
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b1111111011100000,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b1111111100100100,
                    `W_DATA_BITWIDTH'b1111111101101110,
                    `W_DATA_BITWIDTH'b1111111101101100,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111001010001,
                    `W_DATA_BITWIDTH'b1111111101000010,
                    `W_DATA_BITWIDTH'b1111111011111100,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b1111111010111111,
                    `W_DATA_BITWIDTH'b0000000010001010,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b1111111000101010,
                    `W_DATA_BITWIDTH'b0000000100101101,
                    `W_DATA_BITWIDTH'b0000001001100010,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000001010100001,
                    `W_DATA_BITWIDTH'b0000000011001010,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b0000000110001110,
                    `W_DATA_BITWIDTH'b1111111100100001,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b1111111010101101,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000100011010,
                    `W_DATA_BITWIDTH'b1111111100110011,
                    `W_DATA_BITWIDTH'b0000000110101000,
                    `W_DATA_BITWIDTH'b0000000011000000,
                    `W_DATA_BITWIDTH'b0000000111011000,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b0000000111100110,
                    `W_DATA_BITWIDTH'b1111111011111101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000110011101,
                    `W_DATA_BITWIDTH'b1111111101111011,
                    `W_DATA_BITWIDTH'b1111111000111001,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b1111111001001001,
                    `W_DATA_BITWIDTH'b0000000111111000,
                    `W_DATA_BITWIDTH'b1111111001111011,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b1111111011010010,
                    `W_DATA_BITWIDTH'b1111111000011001,
                    `W_DATA_BITWIDTH'b0000000010001010,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111111010000011,
                    `W_DATA_BITWIDTH'b0000000011000110,
                    `W_DATA_BITWIDTH'b1111111001111010,
                    `W_DATA_BITWIDTH'b1111110111011001,
                    `W_DATA_BITWIDTH'b1111111101010001,
                    `W_DATA_BITWIDTH'b1111111001110011,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b0000000101101111,
                    `W_DATA_BITWIDTH'b0000000101011111,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b1111111101110011,
                    `W_DATA_BITWIDTH'b1111111101100010,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111110111100100,
                    `W_DATA_BITWIDTH'b1111111101011111,
                    `W_DATA_BITWIDTH'b0000000011100101,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b1111110110010110,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b0000000110001000,
                    `W_DATA_BITWIDTH'b1111111011101011,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b1111111010001111,
                    `W_DATA_BITWIDTH'b0000000110010101,
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b0000000100000000,
                    `W_DATA_BITWIDTH'b1111111001010000,
                    `W_DATA_BITWIDTH'b0000000011111101,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b0000000010011100,
                    `W_DATA_BITWIDTH'b1111111101111011,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111101001010,
                    `W_DATA_BITWIDTH'b0000000011110101,
                    `W_DATA_BITWIDTH'b0000000100111110,
                    `W_DATA_BITWIDTH'b0000000100011011,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b1111111100110000,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b0000000011101101,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111001111101,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b1111111010011000,
                    `W_DATA_BITWIDTH'b0000000011001001,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000010011010,
                    `W_DATA_BITWIDTH'b0000000100010001,
                    `W_DATA_BITWIDTH'b1111111011011011,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111011011001,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b1111111011100111,
                    `W_DATA_BITWIDTH'b0000000011111110,
                    `W_DATA_BITWIDTH'b0000000100000100,
                    `W_DATA_BITWIDTH'b0000000010100100,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000011110100,
                    `W_DATA_BITWIDTH'b0000000010010000,
                    `W_DATA_BITWIDTH'b0000000010111000,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b0000000010001010,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b0000000010011100,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b1111110111010111,
                    `W_DATA_BITWIDTH'b1111111001100011,
                    `W_DATA_BITWIDTH'b1111110111111111,
                    `W_DATA_BITWIDTH'b1111110110100011,
                    `W_DATA_BITWIDTH'b0000000010110110,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000101110000,
                    `W_DATA_BITWIDTH'b1111111010110011,
                    `W_DATA_BITWIDTH'b1111111101100010,
                    `W_DATA_BITWIDTH'b1111110111001110,
                    `W_DATA_BITWIDTH'b1111110001110100,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111110110011011,
                    `W_DATA_BITWIDTH'b1111111011111001,
                    `W_DATA_BITWIDTH'b1111111011111000,
                    `W_DATA_BITWIDTH'b0000000100011100,
                    `W_DATA_BITWIDTH'b1111111000001101,
                    `W_DATA_BITWIDTH'b0000000100001001,
                    `W_DATA_BITWIDTH'b0000000100111100,
                    `W_DATA_BITWIDTH'b0000000101100110,
                    `W_DATA_BITWIDTH'b0000000101100101,
                    `W_DATA_BITWIDTH'b1111111000010001,
                    `W_DATA_BITWIDTH'b0000000110110101,
                    `W_DATA_BITWIDTH'b0000001000001111,
                    `W_DATA_BITWIDTH'b0000000111011010,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b1111111100001000,
                    `W_DATA_BITWIDTH'b0000000010001110,
                    `W_DATA_BITWIDTH'b1111111011101111,
                    `W_DATA_BITWIDTH'b1111111011001101,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b0000000101010000,
                    `W_DATA_BITWIDTH'b0000000101010000
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
                '{
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111111100100001,
                    `W_DATA_BITWIDTH'b1111111011010011,
                    `W_DATA_BITWIDTH'b1111111010000100,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b1111111011111100,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111111001011101,
                    `W_DATA_BITWIDTH'b1111111100010101,
                    `W_DATA_BITWIDTH'b1111111101010011,
                    `W_DATA_BITWIDTH'b1111111100000110,
                    `W_DATA_BITWIDTH'b1111111001111001,
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b1111111010000001,
                    `W_DATA_BITWIDTH'b0000000011111001,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b1111111100100010,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b0000000010110010,
                    `W_DATA_BITWIDTH'b1111111101100101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b0000000100100110,
                    `W_DATA_BITWIDTH'b0000000010111100,
                    `W_DATA_BITWIDTH'b1111111101100101,
                    `W_DATA_BITWIDTH'b1111111010111001,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b1111111100001100,
                    `W_DATA_BITWIDTH'b1111111010011111,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b0000000011001011,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b0000000011010100,
                    `W_DATA_BITWIDTH'b0000000010000101,
                    `W_DATA_BITWIDTH'b0000000011111010,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b0000000010010001,
                    `W_DATA_BITWIDTH'b0000000011010010,
                    `W_DATA_BITWIDTH'b0000000010010100,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b0000000011111010,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b0000000100111100,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111101000111,
                    `W_DATA_BITWIDTH'b0000000011111010,
                    `W_DATA_BITWIDTH'b0000000011000001,
                    `W_DATA_BITWIDTH'b0000000101000101,
                    `W_DATA_BITWIDTH'b1111111011010000,
                    `W_DATA_BITWIDTH'b1111111001101011,
                    `W_DATA_BITWIDTH'b1111111010100111,
                    `W_DATA_BITWIDTH'b1111111011010001,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000110101011,
                    `W_DATA_BITWIDTH'b0000000011011010,
                    `W_DATA_BITWIDTH'b0000000100010010,
                    `W_DATA_BITWIDTH'b0000000101000000,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000100111011,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b1111111010100001,
                    `W_DATA_BITWIDTH'b0000000101000010,
                    `W_DATA_BITWIDTH'b1111111011101001,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111111010110110,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b1111111010010010,
                    `W_DATA_BITWIDTH'b0000000011111001,
                    `W_DATA_BITWIDTH'b0000000011111001,
                    `W_DATA_BITWIDTH'b1111111001111101,
                    `W_DATA_BITWIDTH'b0000000011101000,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000101011110,
                    `W_DATA_BITWIDTH'b1111110111101100,
                    `W_DATA_BITWIDTH'b0000000110101001,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000100110111,
                    `W_DATA_BITWIDTH'b1111110100110000,
                    `W_DATA_BITWIDTH'b0000000110000111,
                    `W_DATA_BITWIDTH'b1111111011100010,
                    `W_DATA_BITWIDTH'b1111111010000110,
                    `W_DATA_BITWIDTH'b1111111001000001,
                    `W_DATA_BITWIDTH'b1111110100100101,
                    `W_DATA_BITWIDTH'b1111111100101100,
                    `W_DATA_BITWIDTH'b1111111001000111,
                    `W_DATA_BITWIDTH'b0000000011010110,
                    `W_DATA_BITWIDTH'b0000000110101010,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111100000111,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b1111111000001100,
                    `W_DATA_BITWIDTH'b0000000101100111,
                    `W_DATA_BITWIDTH'b0000000111111010,
                    `W_DATA_BITWIDTH'b0000000111010110,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b0000000101001011,
                    `W_DATA_BITWIDTH'b0000000111111000,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b0000000101001000,
                    `W_DATA_BITWIDTH'b1111110100110011,
                    `W_DATA_BITWIDTH'b0000000110100100,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111111011001001,
                    `W_DATA_BITWIDTH'b0000001001110111,
                    `W_DATA_BITWIDTH'b0000001001011010,
                    `W_DATA_BITWIDTH'b0000000011001001,
                    `W_DATA_BITWIDTH'b1111111011101100,
                    `W_DATA_BITWIDTH'b1111111001110110,
                    `W_DATA_BITWIDTH'b0000000010000101,
                    `W_DATA_BITWIDTH'b1111111000101001,
                    `W_DATA_BITWIDTH'b1111111001100101,
                    `W_DATA_BITWIDTH'b0000000101101010,
                    `W_DATA_BITWIDTH'b1111111100111010,
                    `W_DATA_BITWIDTH'b1111111001001101,
                    `W_DATA_BITWIDTH'b1111111101011101,
                    `W_DATA_BITWIDTH'b0000000011010111,
                    `W_DATA_BITWIDTH'b1111110111000101,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111101111111,
                    `W_DATA_BITWIDTH'b1111111100111001,
                    `W_DATA_BITWIDTH'b1111111011100011,
                    `W_DATA_BITWIDTH'b1111111101001001,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011010010,
                    `W_DATA_BITWIDTH'b1111111100100100,
                    `W_DATA_BITWIDTH'b1111111011110000,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b0000000011110010,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111000110011,
                    `W_DATA_BITWIDTH'b0000000101110101,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b0000000010101001,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b1111111100110111,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b0000000100100110,
                    `W_DATA_BITWIDTH'b1111111000010011,
                    `W_DATA_BITWIDTH'b1111111100001001,
                    `W_DATA_BITWIDTH'b1111111101000001,
                    `W_DATA_BITWIDTH'b1111111100011111,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b1111111101101101,
                    `W_DATA_BITWIDTH'b1111111100011010,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000100110011,
                    `W_DATA_BITWIDTH'b0000000100010110,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b1111111100110101,
                    `W_DATA_BITWIDTH'b0000000010101001,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111011000010,
                    `W_DATA_BITWIDTH'b0000000010010101,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b0000000010001000,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b0000000011001010,
                    `W_DATA_BITWIDTH'b1111111101001001,
                    `W_DATA_BITWIDTH'b0000000011010011,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111111100001000,
                    `W_DATA_BITWIDTH'b1111111011010111,
                    `W_DATA_BITWIDTH'b0000000011100001,
                    `W_DATA_BITWIDTH'b0000000101110111,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b1111111011010101,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000010000101,
                    `W_DATA_BITWIDTH'b0000000101110001,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b1111111011000010,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b1111111101110100,
                    `W_DATA_BITWIDTH'b1111111101101110,
                    `W_DATA_BITWIDTH'b1111111101001000,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111101010010,
                    `W_DATA_BITWIDTH'b1111111001110010,
                    `W_DATA_BITWIDTH'b0000000010100000,
                    `W_DATA_BITWIDTH'b1111111100011100,
                    `W_DATA_BITWIDTH'b0000000011110110,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b0000000010101001,
                    `W_DATA_BITWIDTH'b1111111100010110,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b1111111001010000,
                    `W_DATA_BITWIDTH'b1111111011111111,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b1111111011100011,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111010110010,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111111100010111,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000011010010,
                    `W_DATA_BITWIDTH'b0000000110010010,
                    `W_DATA_BITWIDTH'b0000000011110101,
                    `W_DATA_BITWIDTH'b1111111101010110,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000100000100,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b0000000111101000,
                    `W_DATA_BITWIDTH'b0000001000111011,
                    `W_DATA_BITWIDTH'b0000000111010000,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b1111111101100000,
                    `W_DATA_BITWIDTH'b0000000101100011,
                    `W_DATA_BITWIDTH'b1111110110110001,
                    `W_DATA_BITWIDTH'b0000001000011111,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b1111111000011100,
                    `W_DATA_BITWIDTH'b0000000111110101,
                    `W_DATA_BITWIDTH'b1111111100110000,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b1111110110101110,
                    `W_DATA_BITWIDTH'b0000000101000001,
                    `W_DATA_BITWIDTH'b0000000110100011,
                    `W_DATA_BITWIDTH'b0000000100111011,
                    `W_DATA_BITWIDTH'b0000000100001000,
                    `W_DATA_BITWIDTH'b1111110101001010,
                    `W_DATA_BITWIDTH'b1111111000101010,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111100110000,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111110111010001,
                    `W_DATA_BITWIDTH'b1111111101000111,
                    `W_DATA_BITWIDTH'b0000000011110100,
                    `W_DATA_BITWIDTH'b0000000110101110,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000100100111,
                    `W_DATA_BITWIDTH'b1111110111010011,
                    `W_DATA_BITWIDTH'b0000000110101101,
                    `W_DATA_BITWIDTH'b0000000011010110,
                    `W_DATA_BITWIDTH'b0000000101110110,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b0000000011100000,
                    `W_DATA_BITWIDTH'b1111111100111110,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111101101111,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b0000000011011101,
                    `W_DATA_BITWIDTH'b1111111100000011,
                    `W_DATA_BITWIDTH'b1111111011101111,
                    `W_DATA_BITWIDTH'b0000000011011101,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111101010010,
                    `W_DATA_BITWIDTH'b1111111010010101,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b0000000110111111,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b1111111101100000,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b0000001000011001,
                    `W_DATA_BITWIDTH'b1111111010001010,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b1111111100101100,
                    `W_DATA_BITWIDTH'b1111111001110110,
                    `W_DATA_BITWIDTH'b0000000011111101,
                    `W_DATA_BITWIDTH'b0000000100110101,
                    `W_DATA_BITWIDTH'b1111111000111011,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000011010110,
                    `W_DATA_BITWIDTH'b1111111011101111,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111010010011,
                    `W_DATA_BITWIDTH'b1111111100111010,
                    `W_DATA_BITWIDTH'b1111111011111110,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b1111111100001001,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b0000000010011010,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b1111111001110100,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b0000000100110101,
                    `W_DATA_BITWIDTH'b1111111011010100,
                    `W_DATA_BITWIDTH'b0000001000110110,
                    `W_DATA_BITWIDTH'b0000000101100111,
                    `W_DATA_BITWIDTH'b0000000101010011,
                    `W_DATA_BITWIDTH'b1111111001110111,
                    `W_DATA_BITWIDTH'b1111111101000001,
                    `W_DATA_BITWIDTH'b0000000101111101,
                    `W_DATA_BITWIDTH'b1111111010000100,
                    `W_DATA_BITWIDTH'b0000000110011110,
                    `W_DATA_BITWIDTH'b0000000101010101,
                    `W_DATA_BITWIDTH'b0000000100100000,
                    `W_DATA_BITWIDTH'b1111111010100000,
                    `W_DATA_BITWIDTH'b1111110110011101,
                    `W_DATA_BITWIDTH'b1111111101000001,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111100000101,
                    `W_DATA_BITWIDTH'b1111110010111001,
                    `W_DATA_BITWIDTH'b0000001000011100,
                    `W_DATA_BITWIDTH'b0000000010110110,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b1111110010011011,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111110101111011,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b0000000111010110,
                    `W_DATA_BITWIDTH'b1111111100100001,
                    `W_DATA_BITWIDTH'b1111111000100001,
                    `W_DATA_BITWIDTH'b1111111001011001,
                    `W_DATA_BITWIDTH'b1111111010111100,
                    `W_DATA_BITWIDTH'b1111111000101001,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111001000101,
                    `W_DATA_BITWIDTH'b0000000010010010,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111101001000,
                    `W_DATA_BITWIDTH'b1111111101101010,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b1111111011000001,
                    `W_DATA_BITWIDTH'b1111111010110011,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b0000000100011011,
                    `W_DATA_BITWIDTH'b1111111000110110,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111111000010011,
                    `W_DATA_BITWIDTH'b1111111100100101,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b0000000110010110,
                    `W_DATA_BITWIDTH'b0000000010110101,
                    `W_DATA_BITWIDTH'b1111111101001011,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b1111111101100100,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111111100101110,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111111001100011,
                    `W_DATA_BITWIDTH'b0000000110011110,
                    `W_DATA_BITWIDTH'b0000000101110111,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b1111111101101111,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000100101111,
                    `W_DATA_BITWIDTH'b1111111101100001,
                    `W_DATA_BITWIDTH'b0000000101110000,
                    `W_DATA_BITWIDTH'b0000000101010010,
                    `W_DATA_BITWIDTH'b0000000110000111,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000100111110,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b1111111010110101,
                    `W_DATA_BITWIDTH'b1111111101111011,
                    `W_DATA_BITWIDTH'b0000000100010101,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b0000000100001011,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000100000001,
                    `W_DATA_BITWIDTH'b0000000100111111,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111110110110000,
                    `W_DATA_BITWIDTH'b1111111101000011,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b0000000010101010,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b0000000011001101,
                    `W_DATA_BITWIDTH'b0000000100100110,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111111100110010,
                    `W_DATA_BITWIDTH'b0000000010010101,
                    `W_DATA_BITWIDTH'b0000000101010110,
                    `W_DATA_BITWIDTH'b0000000011011000,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b0000000011100010,
                    `W_DATA_BITWIDTH'b1111111101110100,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b0000000100100010,
                    `W_DATA_BITWIDTH'b0000000011010111,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111100000101,
                    `W_DATA_BITWIDTH'b1111110110010000,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b1111111011111011,
                    `W_DATA_BITWIDTH'b1111111011100001,
                    `W_DATA_BITWIDTH'b0000000101011000,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000011011000,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111110110101100,
                    `W_DATA_BITWIDTH'b1111111100010110,
                    `W_DATA_BITWIDTH'b1111111100001100,
                    `W_DATA_BITWIDTH'b1111111100100101,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b1111111010001110,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b1111111000010010,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b1111111010001110,
                    `W_DATA_BITWIDTH'b1111111010110101,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111100000101,
                    `W_DATA_BITWIDTH'b1111111000000110,
                    `W_DATA_BITWIDTH'b1111111101100010,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b0000000100100010,
                    `W_DATA_BITWIDTH'b0000000110000001,
                    `W_DATA_BITWIDTH'b0000000100000000,
                    `W_DATA_BITWIDTH'b0000001001000010,
                    `W_DATA_BITWIDTH'b0000001001000010
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000010100010,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b1111111101100100,
                    `W_DATA_BITWIDTH'b0000000011010001,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b0000000011010100,
                    `W_DATA_BITWIDTH'b1111111011110100,
                    `W_DATA_BITWIDTH'b1111111010010100,
                    `W_DATA_BITWIDTH'b0000000010010010,
                    `W_DATA_BITWIDTH'b1111111001110100,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b1111111100111010,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b0000000100110101,
                    `W_DATA_BITWIDTH'b1111111011111001,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b0000000101001111,
                    `W_DATA_BITWIDTH'b1111111101011000,
                    `W_DATA_BITWIDTH'b0000000100000010,
                    `W_DATA_BITWIDTH'b1111111100101010,
                    `W_DATA_BITWIDTH'b1111111011001011,
                    `W_DATA_BITWIDTH'b1111111100100110,
                    `W_DATA_BITWIDTH'b0000000010010000,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b1111111011111100,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b0000000100101100,
                    `W_DATA_BITWIDTH'b0000000010101010,
                    `W_DATA_BITWIDTH'b0000000100101011,
                    `W_DATA_BITWIDTH'b1111111101010011,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b1111111010110010,
                    `W_DATA_BITWIDTH'b1111111010000100,
                    `W_DATA_BITWIDTH'b1111111101000110,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b0000000101000111,
                    `W_DATA_BITWIDTH'b0000001000110101,
                    `W_DATA_BITWIDTH'b1111111010010101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011111111,
                    `W_DATA_BITWIDTH'b0000000011100110,
                    `W_DATA_BITWIDTH'b1111111010000101,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111101110001,
                    `W_DATA_BITWIDTH'b0000000011100111,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000000011011010,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b0000000011101100,
                    `W_DATA_BITWIDTH'b0000000100011001,
                    `W_DATA_BITWIDTH'b1111111000101110,
                    `W_DATA_BITWIDTH'b0000000111111110,
                    `W_DATA_BITWIDTH'b1111111001111000,
                    `W_DATA_BITWIDTH'b1111111100110011,
                    `W_DATA_BITWIDTH'b1111111000101101,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b1111110111100011,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b0000001011111010,
                    `W_DATA_BITWIDTH'b0000000100011000,
                    `W_DATA_BITWIDTH'b0000000110000001,
                    `W_DATA_BITWIDTH'b1111111011100101,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b1111110111100100,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b0000000101101110,
                    `W_DATA_BITWIDTH'b0000000011111110,
                    `W_DATA_BITWIDTH'b0000001000101110,
                    `W_DATA_BITWIDTH'b1111111000011001,
                    `W_DATA_BITWIDTH'b0000000100000001,
                    `W_DATA_BITWIDTH'b0000000101010111,
                    `W_DATA_BITWIDTH'b1111111001001100,
                    `W_DATA_BITWIDTH'b1111111011111101,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000110101010,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b1111111001011101,
                    `W_DATA_BITWIDTH'b1111111100001100,
                    `W_DATA_BITWIDTH'b0000000010101010,
                    `W_DATA_BITWIDTH'b1111110110110001,
                    `W_DATA_BITWIDTH'b1111111101101101,
                    `W_DATA_BITWIDTH'b1111110110111000,
                    `W_DATA_BITWIDTH'b0000001010000111,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b0000000100100111,
                    `W_DATA_BITWIDTH'b0000000100000001,
                    `W_DATA_BITWIDTH'b1111110110111110,
                    `W_DATA_BITWIDTH'b0000000110101001,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b1111110100100011,
                    `W_DATA_BITWIDTH'b0000000011101100,
                    `W_DATA_BITWIDTH'b1111111000000111,
                    `W_DATA_BITWIDTH'b1111111100001011,
                    `W_DATA_BITWIDTH'b1111111011010000,
                    `W_DATA_BITWIDTH'b1111111001000101,
                    `W_DATA_BITWIDTH'b1111111101011111,
                    `W_DATA_BITWIDTH'b1111110110100000,
                    `W_DATA_BITWIDTH'b1111111001111111,
                    `W_DATA_BITWIDTH'b0000000101101110,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b1111111001111010,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b0000000100010011,
                    `W_DATA_BITWIDTH'b1111111011010001,
                    `W_DATA_BITWIDTH'b0000000101010111,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b1111111100010111,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111100111101,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b0000000011111111,
                    `W_DATA_BITWIDTH'b0000000101011001,
                    `W_DATA_BITWIDTH'b0000000011010100,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b1111111101011001,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b1111111010001001,
                    `W_DATA_BITWIDTH'b0000000100000111,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b0000000010011001,
                    `W_DATA_BITWIDTH'b1111111100010011,
                    `W_DATA_BITWIDTH'b1111111001111111,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111011100000,
                    `W_DATA_BITWIDTH'b0000000101111010,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111001111010,
                    `W_DATA_BITWIDTH'b0000000011101100,
                    `W_DATA_BITWIDTH'b1111111011001000,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b1111111001100100,
                    `W_DATA_BITWIDTH'b0000000100100000,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b1111111011110010,
                    `W_DATA_BITWIDTH'b1111110111010100,
                    `W_DATA_BITWIDTH'b1111111011101101,
                    `W_DATA_BITWIDTH'b1111111011001010,
                    `W_DATA_BITWIDTH'b1111111001101101,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000010011101,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000100111000,
                    `W_DATA_BITWIDTH'b1111111001111100,
                    `W_DATA_BITWIDTH'b1111111101010011,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000011011111,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b1111110111101111,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b1111111100111101,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b0000000100100011,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111110110101010,
                    `W_DATA_BITWIDTH'b1111111010011000,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111001111101,
                    `W_DATA_BITWIDTH'b1111111011011101,
                    `W_DATA_BITWIDTH'b1111111010101100,
                    `W_DATA_BITWIDTH'b0000000010001000,
                    `W_DATA_BITWIDTH'b1111111000110010,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b1111111011001001,
                    `W_DATA_BITWIDTH'b0000000011111000,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b1111111011011011,
                    `W_DATA_BITWIDTH'b1111111011000010,
                    `W_DATA_BITWIDTH'b1111111010111111,
                    `W_DATA_BITWIDTH'b1111111011101100,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111010011101,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b0000000011000001,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b1111111101001110,
                    `W_DATA_BITWIDTH'b1111111010110011,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b1111111010101000,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b1111111000011101,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b0000000101100101,
                    `W_DATA_BITWIDTH'b0000000101000110,
                    `W_DATA_BITWIDTH'b1111111011011100,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111000110101,
                    `W_DATA_BITWIDTH'b0000000100100111,
                    `W_DATA_BITWIDTH'b1111110010101100,
                    `W_DATA_BITWIDTH'b1111110101111001,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b1111111010010111,
                    `W_DATA_BITWIDTH'b1111111001100101,
                    `W_DATA_BITWIDTH'b0000000101010110,
                    `W_DATA_BITWIDTH'b0000000010011001,
                    `W_DATA_BITWIDTH'b0000001010001010,
                    `W_DATA_BITWIDTH'b1111111000111101,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b1111111001000111,
                    `W_DATA_BITWIDTH'b1111111010100111,
                    `W_DATA_BITWIDTH'b1111111000110000,
                    `W_DATA_BITWIDTH'b1111111000101011,
                    `W_DATA_BITWIDTH'b0000000100100000,
                    `W_DATA_BITWIDTH'b0000000011011011,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b0000000111001010,
                    `W_DATA_BITWIDTH'b0000000101001000,
                    `W_DATA_BITWIDTH'b1111111001011001,
                    `W_DATA_BITWIDTH'b0000000101011010,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111111101111110,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b0000000011110000,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b1111111100111101,
                    `W_DATA_BITWIDTH'b0000000100001100,
                    `W_DATA_BITWIDTH'b0000000101000100,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000011001010,
                    `W_DATA_BITWIDTH'b1111111011110010,
                    `W_DATA_BITWIDTH'b1111111011101011,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000100001011,
                    `W_DATA_BITWIDTH'b0000000011110000,
                    `W_DATA_BITWIDTH'b1111111011000011,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111111101111000,
                    `W_DATA_BITWIDTH'b0000000101010111,
                    `W_DATA_BITWIDTH'b0000000010010001,
                    `W_DATA_BITWIDTH'b1111111101011110,
                    `W_DATA_BITWIDTH'b0000000110110001,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b0000001000001001,
                    `W_DATA_BITWIDTH'b0000000010011010,
                    `W_DATA_BITWIDTH'b0000000100011010,
                    `W_DATA_BITWIDTH'b0000000110010110,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b0000000110111000,
                    `W_DATA_BITWIDTH'b0000000011111101,
                    `W_DATA_BITWIDTH'b1111111001011110,
                    `W_DATA_BITWIDTH'b0000000011111011,
                    `W_DATA_BITWIDTH'b1111111100010100,
                    `W_DATA_BITWIDTH'b0000000011101101,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b1111111100111001,
                    `W_DATA_BITWIDTH'b0000000010100000,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b1111110111110110,
                    `W_DATA_BITWIDTH'b0000000101110100,
                    `W_DATA_BITWIDTH'b0000000110001101,
                    `W_DATA_BITWIDTH'b1111111001110000,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b0000000010001110,
                    `W_DATA_BITWIDTH'b0000000101110011,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b1111110101111011,
                    `W_DATA_BITWIDTH'b0000001001101010,
                    `W_DATA_BITWIDTH'b0000000100110000,
                    `W_DATA_BITWIDTH'b1111110001100010,
                    `W_DATA_BITWIDTH'b0000001001110100,
                    `W_DATA_BITWIDTH'b0000000111000100,
                    `W_DATA_BITWIDTH'b1111111011110111,
                    `W_DATA_BITWIDTH'b1111110110100111,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b1111111000001000,
                    `W_DATA_BITWIDTH'b1111111101001000,
                    `W_DATA_BITWIDTH'b0000000110011101,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b1111110100100100,
                    `W_DATA_BITWIDTH'b0000000101000100,
                    `W_DATA_BITWIDTH'b0000000110101011,
                    `W_DATA_BITWIDTH'b1111111010111010,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b1111111101011100,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b0000000101100010,
                    `W_DATA_BITWIDTH'b1111111000011100,
                    `W_DATA_BITWIDTH'b0000000011001011,
                    `W_DATA_BITWIDTH'b1111111100000011,
                    `W_DATA_BITWIDTH'b1111111011010111,
                    `W_DATA_BITWIDTH'b0000000101111110,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111110011111000,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b0000000010100101,
                    `W_DATA_BITWIDTH'b1111111011100011,
                    `W_DATA_BITWIDTH'b1111111001001100,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b1111111001110010,
                    `W_DATA_BITWIDTH'b1111111101110100,
                    `W_DATA_BITWIDTH'b0000000101101000,
                    `W_DATA_BITWIDTH'b1111111001101100,
                    `W_DATA_BITWIDTH'b1111111010110000,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b0000000011111011,
                    `W_DATA_BITWIDTH'b1111111010010100,
                    `W_DATA_BITWIDTH'b0000000101010000,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b1111111000101000,
                    `W_DATA_BITWIDTH'b1111111100111100,
                    `W_DATA_BITWIDTH'b0000000101001000,
                    `W_DATA_BITWIDTH'b0000000110000010,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b0000000010110101,
                    `W_DATA_BITWIDTH'b1111111001011100,
                    `W_DATA_BITWIDTH'b0000000011001110,
                    `W_DATA_BITWIDTH'b1111111100010101,
                    `W_DATA_BITWIDTH'b1111111101001101,
                    `W_DATA_BITWIDTH'b1111111011011111,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b1111111010101110,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b1111111100100010,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b0000000100001000,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000101000101,
                    `W_DATA_BITWIDTH'b0000000011000001,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b1111111011111111,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b0000000010111100,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b0000000100101011,
                    `W_DATA_BITWIDTH'b0000000101101101,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b1111110101001100,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111011111101,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b0000000100101111,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b0000000010001110,
                    `W_DATA_BITWIDTH'b1111111101100001,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b0000000100000111,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b1111111011000001,
                    `W_DATA_BITWIDTH'b1111111001100000,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b1111110110000111,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b1111111010011101,
                    `W_DATA_BITWIDTH'b0000000101000110,
                    `W_DATA_BITWIDTH'b0000000101100011,
                    `W_DATA_BITWIDTH'b0000000010100101,
                    `W_DATA_BITWIDTH'b0000000101011011,
                    `W_DATA_BITWIDTH'b1111111100011111,
                    `W_DATA_BITWIDTH'b1111111001100010,
                    `W_DATA_BITWIDTH'b0000000100011000,
                    `W_DATA_BITWIDTH'b0000000100010011,
                    `W_DATA_BITWIDTH'b1111111101110011,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b0000000100111011,
                    `W_DATA_BITWIDTH'b1111111010001011,
                    `W_DATA_BITWIDTH'b1111111100000111,
                    `W_DATA_BITWIDTH'b0000001001000101,
                    `W_DATA_BITWIDTH'b1111111101001111,
                    `W_DATA_BITWIDTH'b1111111010010110,
                    `W_DATA_BITWIDTH'b0000001000111001,
                    `W_DATA_BITWIDTH'b0000000111110000,
                    `W_DATA_BITWIDTH'b1111111101101001,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b1111111011001000,
                    `W_DATA_BITWIDTH'b0000000011011011,
                    `W_DATA_BITWIDTH'b1111110110110101,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b0000000100000110,
                    `W_DATA_BITWIDTH'b0000001000000111,
                    `W_DATA_BITWIDTH'b0000000100111100,
                    `W_DATA_BITWIDTH'b0000000100111100
                };

            // w_c_idx
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
                '{
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
                '{
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
                '{
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
                '{
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01110
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
                '{
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01110
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
                '{
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01110
                };

            // w_r_idx
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };

            // w_k_idx
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };

            // w_pos_ptr
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00000000000,
                    `W_POS_PTR_BITWIDTH'b00000000010,
                    `W_POS_PTR_BITWIDTH'b00000000100,
                    `W_POS_PTR_BITWIDTH'b00000000110,
                    `W_POS_PTR_BITWIDTH'b00000001000,
                    `W_POS_PTR_BITWIDTH'b00000001010,
                    `W_POS_PTR_BITWIDTH'b00000001101,
                    `W_POS_PTR_BITWIDTH'b00000010000,
                    `W_POS_PTR_BITWIDTH'b00000010011,
                    `W_POS_PTR_BITWIDTH'b00000010110,
                    `W_POS_PTR_BITWIDTH'b00000011001,
                    `W_POS_PTR_BITWIDTH'b00000011100,
                    `W_POS_PTR_BITWIDTH'b00000011110,
                    `W_POS_PTR_BITWIDTH'b00000100000,
                    `W_POS_PTR_BITWIDTH'b00000100011,
                    `W_POS_PTR_BITWIDTH'b00000100110,
                    `W_POS_PTR_BITWIDTH'b00000101001,
                    `W_POS_PTR_BITWIDTH'b00000101100,
                    `W_POS_PTR_BITWIDTH'b00000101110,
                    `W_POS_PTR_BITWIDTH'b00000110000,
                    `W_POS_PTR_BITWIDTH'b00000110011,
                    `W_POS_PTR_BITWIDTH'b00000110101,
                    `W_POS_PTR_BITWIDTH'b00000111000,
                    `W_POS_PTR_BITWIDTH'b00000111010,
                    `W_POS_PTR_BITWIDTH'b00000111100,
                    `W_POS_PTR_BITWIDTH'b00000111111,
                    `W_POS_PTR_BITWIDTH'b00001000010,
                    `W_POS_PTR_BITWIDTH'b00001000100,
                    `W_POS_PTR_BITWIDTH'b00001000111,
                    `W_POS_PTR_BITWIDTH'b00001001010,
                    `W_POS_PTR_BITWIDTH'b00001001101,
                    `W_POS_PTR_BITWIDTH'b00001001110,
                    `W_POS_PTR_BITWIDTH'b00001010000,
                    `W_POS_PTR_BITWIDTH'b00001010010,
                    `W_POS_PTR_BITWIDTH'b00001010101,
                    `W_POS_PTR_BITWIDTH'b00001011000,
                    `W_POS_PTR_BITWIDTH'b00001011011,
                    `W_POS_PTR_BITWIDTH'b00001011110,
                    `W_POS_PTR_BITWIDTH'b00001100001,
                    `W_POS_PTR_BITWIDTH'b00001100100,
                    `W_POS_PTR_BITWIDTH'b00001100110,
                    `W_POS_PTR_BITWIDTH'b00001101000,
                    `W_POS_PTR_BITWIDTH'b00001101011,
                    `W_POS_PTR_BITWIDTH'b00001101101,
                    `W_POS_PTR_BITWIDTH'b00001110000,
                    `W_POS_PTR_BITWIDTH'b00001110010,
                    `W_POS_PTR_BITWIDTH'b00001110101,
                    `W_POS_PTR_BITWIDTH'b00001110101
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00001111011,
                    `W_POS_PTR_BITWIDTH'b00001111101,
                    `W_POS_PTR_BITWIDTH'b00001111111,
                    `W_POS_PTR_BITWIDTH'b00010000010,
                    `W_POS_PTR_BITWIDTH'b00010000101,
                    `W_POS_PTR_BITWIDTH'b00010001000,
                    `W_POS_PTR_BITWIDTH'b00010001011,
                    `W_POS_PTR_BITWIDTH'b00010001110,
                    `W_POS_PTR_BITWIDTH'b00010010001,
                    `W_POS_PTR_BITWIDTH'b00010010100,
                    `W_POS_PTR_BITWIDTH'b00010010111,
                    `W_POS_PTR_BITWIDTH'b00010011001,
                    `W_POS_PTR_BITWIDTH'b00010011100,
                    `W_POS_PTR_BITWIDTH'b00010011111,
                    `W_POS_PTR_BITWIDTH'b00010100010,
                    `W_POS_PTR_BITWIDTH'b00010100101,
                    `W_POS_PTR_BITWIDTH'b00010101000,
                    `W_POS_PTR_BITWIDTH'b00010101011,
                    `W_POS_PTR_BITWIDTH'b00010101110,
                    `W_POS_PTR_BITWIDTH'b00010110000,
                    `W_POS_PTR_BITWIDTH'b00010110010,
                    `W_POS_PTR_BITWIDTH'b00010110101,
                    `W_POS_PTR_BITWIDTH'b00010111000,
                    `W_POS_PTR_BITWIDTH'b00010111010,
                    `W_POS_PTR_BITWIDTH'b00010111101,
                    `W_POS_PTR_BITWIDTH'b00011000000,
                    `W_POS_PTR_BITWIDTH'b00011000011,
                    `W_POS_PTR_BITWIDTH'b00011000110,
                    `W_POS_PTR_BITWIDTH'b00011001001,
                    `W_POS_PTR_BITWIDTH'b00011001100,
                    `W_POS_PTR_BITWIDTH'b00011001110,
                    `W_POS_PTR_BITWIDTH'b00011010000,
                    `W_POS_PTR_BITWIDTH'b00011010010,
                    `W_POS_PTR_BITWIDTH'b00011010011,
                    `W_POS_PTR_BITWIDTH'b00011010110,
                    `W_POS_PTR_BITWIDTH'b00011011001,
                    `W_POS_PTR_BITWIDTH'b00011011100,
                    `W_POS_PTR_BITWIDTH'b00011011111,
                    `W_POS_PTR_BITWIDTH'b00011100010,
                    `W_POS_PTR_BITWIDTH'b00011100101,
                    `W_POS_PTR_BITWIDTH'b00011101000,
                    `W_POS_PTR_BITWIDTH'b00011101011,
                    `W_POS_PTR_BITWIDTH'b00011101110,
                    `W_POS_PTR_BITWIDTH'b00011110000,
                    `W_POS_PTR_BITWIDTH'b00011110010,
                    `W_POS_PTR_BITWIDTH'b00011110101,
                    `W_POS_PTR_BITWIDTH'b00011111000,
                    `W_POS_PTR_BITWIDTH'b00011111000
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00011111101,
                    `W_POS_PTR_BITWIDTH'b00100000000,
                    `W_POS_PTR_BITWIDTH'b00100000010,
                    `W_POS_PTR_BITWIDTH'b00100000101,
                    `W_POS_PTR_BITWIDTH'b00100001000,
                    `W_POS_PTR_BITWIDTH'b00100001001,
                    `W_POS_PTR_BITWIDTH'b00100001100,
                    `W_POS_PTR_BITWIDTH'b00100001111,
                    `W_POS_PTR_BITWIDTH'b00100010010,
                    `W_POS_PTR_BITWIDTH'b00100010101,
                    `W_POS_PTR_BITWIDTH'b00100011000,
                    `W_POS_PTR_BITWIDTH'b00100011011,
                    `W_POS_PTR_BITWIDTH'b00100011110,
                    `W_POS_PTR_BITWIDTH'b00100100000,
                    `W_POS_PTR_BITWIDTH'b00100100011,
                    `W_POS_PTR_BITWIDTH'b00100100110,
                    `W_POS_PTR_BITWIDTH'b00100101000,
                    `W_POS_PTR_BITWIDTH'b00100101011,
                    `W_POS_PTR_BITWIDTH'b00100101110,
                    `W_POS_PTR_BITWIDTH'b00100110000,
                    `W_POS_PTR_BITWIDTH'b00100110011,
                    `W_POS_PTR_BITWIDTH'b00100110110,
                    `W_POS_PTR_BITWIDTH'b00100111000,
                    `W_POS_PTR_BITWIDTH'b00100111010,
                    `W_POS_PTR_BITWIDTH'b00100111101,
                    `W_POS_PTR_BITWIDTH'b00101000000,
                    `W_POS_PTR_BITWIDTH'b00101000011,
                    `W_POS_PTR_BITWIDTH'b00101000110,
                    `W_POS_PTR_BITWIDTH'b00101001001,
                    `W_POS_PTR_BITWIDTH'b00101001100,
                    `W_POS_PTR_BITWIDTH'b00101001111,
                    `W_POS_PTR_BITWIDTH'b00101010000,
                    `W_POS_PTR_BITWIDTH'b00101010001,
                    `W_POS_PTR_BITWIDTH'b00101010010,
                    `W_POS_PTR_BITWIDTH'b00101010100,
                    `W_POS_PTR_BITWIDTH'b00101010111,
                    `W_POS_PTR_BITWIDTH'b00101011010,
                    `W_POS_PTR_BITWIDTH'b00101011101,
                    `W_POS_PTR_BITWIDTH'b00101011111,
                    `W_POS_PTR_BITWIDTH'b00101100010,
                    `W_POS_PTR_BITWIDTH'b00101100100,
                    `W_POS_PTR_BITWIDTH'b00101100111,
                    `W_POS_PTR_BITWIDTH'b00101101010,
                    `W_POS_PTR_BITWIDTH'b00101101100,
                    `W_POS_PTR_BITWIDTH'b00101101110,
                    `W_POS_PTR_BITWIDTH'b00101110001,
                    `W_POS_PTR_BITWIDTH'b00101110100,
                    `W_POS_PTR_BITWIDTH'b00101110100
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00000000000,
                    `W_POS_PTR_BITWIDTH'b00000001010,
                    `W_POS_PTR_BITWIDTH'b00000010001,
                    `W_POS_PTR_BITWIDTH'b00000011001,
                    `W_POS_PTR_BITWIDTH'b00000011111,
                    `W_POS_PTR_BITWIDTH'b00000101001,
                    `W_POS_PTR_BITWIDTH'b00000110001,
                    `W_POS_PTR_BITWIDTH'b00000111001,
                    `W_POS_PTR_BITWIDTH'b00001000101,
                    `W_POS_PTR_BITWIDTH'b00001010001,
                    `W_POS_PTR_BITWIDTH'b00001011110,
                    `W_POS_PTR_BITWIDTH'b00001100110,
                    `W_POS_PTR_BITWIDTH'b00001110100,
                    `W_POS_PTR_BITWIDTH'b00001111111,
                    `W_POS_PTR_BITWIDTH'b00010001001,
                    `W_POS_PTR_BITWIDTH'b00010010100,
                    `W_POS_PTR_BITWIDTH'b00010011011,
                    `W_POS_PTR_BITWIDTH'b00010100101,
                    `W_POS_PTR_BITWIDTH'b00010101110,
                    `W_POS_PTR_BITWIDTH'b00010110101,
                    `W_POS_PTR_BITWIDTH'b00010111110,
                    `W_POS_PTR_BITWIDTH'b00011000100,
                    `W_POS_PTR_BITWIDTH'b00011001101,
                    `W_POS_PTR_BITWIDTH'b00011010110,
                    `W_POS_PTR_BITWIDTH'b00011100000,
                    `W_POS_PTR_BITWIDTH'b00011101011,
                    `W_POS_PTR_BITWIDTH'b00011111000,
                    `W_POS_PTR_BITWIDTH'b00100000110,
                    `W_POS_PTR_BITWIDTH'b00100010000,
                    `W_POS_PTR_BITWIDTH'b00100011001,
                    `W_POS_PTR_BITWIDTH'b00100011110,
                    `W_POS_PTR_BITWIDTH'b00100101001,
                    `W_POS_PTR_BITWIDTH'b00100110111,
                    `W_POS_PTR_BITWIDTH'b00101000000,
                    `W_POS_PTR_BITWIDTH'b00101001010,
                    `W_POS_PTR_BITWIDTH'b00101010100,
                    `W_POS_PTR_BITWIDTH'b00101100001,
                    `W_POS_PTR_BITWIDTH'b00101101101,
                    `W_POS_PTR_BITWIDTH'b00101110111,
                    `W_POS_PTR_BITWIDTH'b00110000011,
                    `W_POS_PTR_BITWIDTH'b00110001101,
                    `W_POS_PTR_BITWIDTH'b00110010110,
                    `W_POS_PTR_BITWIDTH'b00110011110,
                    `W_POS_PTR_BITWIDTH'b00110100101,
                    `W_POS_PTR_BITWIDTH'b00110101111,
                    `W_POS_PTR_BITWIDTH'b00110110110,
                    `W_POS_PTR_BITWIDTH'b00111000011,
                    `W_POS_PTR_BITWIDTH'b00111000011
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00111011010,
                    `W_POS_PTR_BITWIDTH'b00111100100,
                    `W_POS_PTR_BITWIDTH'b00111101110,
                    `W_POS_PTR_BITWIDTH'b00111110111,
                    `W_POS_PTR_BITWIDTH'b01000000000,
                    `W_POS_PTR_BITWIDTH'b01000001000,
                    `W_POS_PTR_BITWIDTH'b01000001110,
                    `W_POS_PTR_BITWIDTH'b01000011000,
                    `W_POS_PTR_BITWIDTH'b01000011110,
                    `W_POS_PTR_BITWIDTH'b01000101010,
                    `W_POS_PTR_BITWIDTH'b01000110101,
                    `W_POS_PTR_BITWIDTH'b01001000010,
                    `W_POS_PTR_BITWIDTH'b01001001111,
                    `W_POS_PTR_BITWIDTH'b01001011100,
                    `W_POS_PTR_BITWIDTH'b01001100001,
                    `W_POS_PTR_BITWIDTH'b01001101011,
                    `W_POS_PTR_BITWIDTH'b01001110100,
                    `W_POS_PTR_BITWIDTH'b01001111100,
                    `W_POS_PTR_BITWIDTH'b01010000100,
                    `W_POS_PTR_BITWIDTH'b01010001111,
                    `W_POS_PTR_BITWIDTH'b01010010111,
                    `W_POS_PTR_BITWIDTH'b01010011110,
                    `W_POS_PTR_BITWIDTH'b01010101010,
                    `W_POS_PTR_BITWIDTH'b01010110010,
                    `W_POS_PTR_BITWIDTH'b01010111110,
                    `W_POS_PTR_BITWIDTH'b01011001000,
                    `W_POS_PTR_BITWIDTH'b01011010101,
                    `W_POS_PTR_BITWIDTH'b01011100010,
                    `W_POS_PTR_BITWIDTH'b01011100111,
                    `W_POS_PTR_BITWIDTH'b01011101111,
                    `W_POS_PTR_BITWIDTH'b01011110100,
                    `W_POS_PTR_BITWIDTH'b01100000000,
                    `W_POS_PTR_BITWIDTH'b01100001000,
                    `W_POS_PTR_BITWIDTH'b01100010001,
                    `W_POS_PTR_BITWIDTH'b01100011011,
                    `W_POS_PTR_BITWIDTH'b01100100101,
                    `W_POS_PTR_BITWIDTH'b01100110100,
                    `W_POS_PTR_BITWIDTH'b01100111111,
                    `W_POS_PTR_BITWIDTH'b01101001000,
                    `W_POS_PTR_BITWIDTH'b01101010011,
                    `W_POS_PTR_BITWIDTH'b01101011111,
                    `W_POS_PTR_BITWIDTH'b01101100111,
                    `W_POS_PTR_BITWIDTH'b01101101101,
                    `W_POS_PTR_BITWIDTH'b01101110111,
                    `W_POS_PTR_BITWIDTH'b01101111110,
                    `W_POS_PTR_BITWIDTH'b01110000101,
                    `W_POS_PTR_BITWIDTH'b01110010001,
                    `W_POS_PTR_BITWIDTH'b01110010001
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b01110100110,
                    `W_POS_PTR_BITWIDTH'b01110101100,
                    `W_POS_PTR_BITWIDTH'b01110110011,
                    `W_POS_PTR_BITWIDTH'b01110111011,
                    `W_POS_PTR_BITWIDTH'b01111000011,
                    `W_POS_PTR_BITWIDTH'b01111001011,
                    `W_POS_PTR_BITWIDTH'b01111010010,
                    `W_POS_PTR_BITWIDTH'b01111011110,
                    `W_POS_PTR_BITWIDTH'b01111100111,
                    `W_POS_PTR_BITWIDTH'b01111110001,
                    `W_POS_PTR_BITWIDTH'b01111111101,
                    `W_POS_PTR_BITWIDTH'b10000001001,
                    `W_POS_PTR_BITWIDTH'b10000010101,
                    `W_POS_PTR_BITWIDTH'b10000011111,
                    `W_POS_PTR_BITWIDTH'b10000100111,
                    `W_POS_PTR_BITWIDTH'b10000110100,
                    `W_POS_PTR_BITWIDTH'b10000111100,
                    `W_POS_PTR_BITWIDTH'b10001000110,
                    `W_POS_PTR_BITWIDTH'b10001001110,
                    `W_POS_PTR_BITWIDTH'b10001010100,
                    `W_POS_PTR_BITWIDTH'b10001100001,
                    `W_POS_PTR_BITWIDTH'b10001101100,
                    `W_POS_PTR_BITWIDTH'b10001110111,
                    `W_POS_PTR_BITWIDTH'b10010000000,
                    `W_POS_PTR_BITWIDTH'b10010000110,
                    `W_POS_PTR_BITWIDTH'b10010010001,
                    `W_POS_PTR_BITWIDTH'b10010011011,
                    `W_POS_PTR_BITWIDTH'b10010101001,
                    `W_POS_PTR_BITWIDTH'b10010110010,
                    `W_POS_PTR_BITWIDTH'b10010111000,
                    `W_POS_PTR_BITWIDTH'b10011000000,
                    `W_POS_PTR_BITWIDTH'b10011001011,
                    `W_POS_PTR_BITWIDTH'b10011010100,
                    `W_POS_PTR_BITWIDTH'b10011011100,
                    `W_POS_PTR_BITWIDTH'b10011101100,
                    `W_POS_PTR_BITWIDTH'b10011110111,
                    `W_POS_PTR_BITWIDTH'b10100000011,
                    `W_POS_PTR_BITWIDTH'b10100001100,
                    `W_POS_PTR_BITWIDTH'b10100010101,
                    `W_POS_PTR_BITWIDTH'b10100011110,
                    `W_POS_PTR_BITWIDTH'b10100100011,
                    `W_POS_PTR_BITWIDTH'b10100101100,
                    `W_POS_PTR_BITWIDTH'b10100110100,
                    `W_POS_PTR_BITWIDTH'b10100111011,
                    `W_POS_PTR_BITWIDTH'b10100111111,
                    `W_POS_PTR_BITWIDTH'b10101000001,
                    `W_POS_PTR_BITWIDTH'b10101001101,
                    `W_POS_PTR_BITWIDTH'b10101001101
                };

        // ----- State ----------
            localparam S_IDLE           = 0;
            localparam S_CAMERA         = 1;

            localparam S_PUT_W_1        = 2;
            localparam S_CONV_1         = 3;
            localparam S_REDUCE_1       = 4;
            localparam S_TOOABUFFER_1   = 5;  // put to OA
            localparam S_COMPRESS_1     = 6;  // put to IA

            localparam S_PUT_W_2        = 7;
            localparam S_CONV_2         = 8;
            localparam S_REDUCE_2       = 9;
            localparam S_TOOABUFFER_2   = 10; // put to OA

            localparam S_MAXPOOL        = 11;
            localparam S_LINEAR         = 12;
            localparam S_OUT            = 13; 

        // ----- PE -----------------
            localparam  logic  PEs_FINISH [0:`PE_ROW-1][0:`PE_COL-1] = 
            '{
                '{1, 1, 1},
                '{1, 1, 1},
                '{1, 1, 1},
                '{1, 1, 1},
                '{1, 1, 1},
                '{1, 1, 1},
                '{1, 1, 1}
            };

            localparam logic  [1:0]                     w_s     [0:`PE_COL-1] = '{0, 1, 2};


            localparam logic  [$clog2(`W_C_LENGTH):0] w_len_1 [0:`PE_COL-1] =
            '{
                `W_C_LENGTH_L1_S0, `W_C_LENGTH_L1_S1, `W_C_LENGTH_L1_S2
            };
            localparam logic  [$clog2(`W_C_LENGTH):0] w_len_2 [0:`PE_COL-1] =
            '{
                `W_C_LENGTH_L2_S0, `W_C_LENGTH_L2_S1, `W_C_LENGTH_L2_S2
            };


            localparam logic  [$clog2(`W_C_LENGTH):0] w_iters_1 [0:`PE_COL-1] =
            '{
                (`W_C_LENGTH_L1_S0 >> 5), (`W_C_LENGTH_L1_S1 >> 5), (`W_C_LENGTH_L1_S2 >>5)
            };
            localparam logic  [$clog2(`W_C_LENGTH):0] w_iters_2 [0:`PE_COL-1] =
            '{
                (`W_C_LENGTH_L2_S0 >> 5), (`W_C_LENGTH_L2_S1 >> 5), (`W_C_LENGTH_L2_S2 >>5)
            };


              


    // ========================== Output Logic ============================================
        logic  [3:0] o_random_out_n;

    // ========================== Logic (Wire) =============================================
        // ----------------------- For PE ------- unfinished------------------------
            
            // IA bundle
            logic        [$clog2(`IA_ROW):0]     i_ia_h      [0:`PE_ROW-1];
            logic        [$clog2(`IA_COL):0]     i_ia_w      [0:`PE_ROW-1];
            logic signed [`IA_DATA_BITWIDTH-1:0]   i_ia_data   [0:`PE_ROW-1][0:`IA_CHANNEL-1];
            logic        [`IA_C_BITWIDTH-1:0]      i_ia_c_idx  [0:`PE_ROW-1][0:`IA_CHANNEL-1];
            logic        [$clog2(`IA_CHANNEL):0] i_ia_iters  [0:`PE_ROW-1];
            logic        [$clog2(`IA_CHANNEL):0] i_ia_len    [0:`PE_ROW-1];
        
            // W bundle
            logic signed [`W_DATA_BITWIDTH-1:0]    i_w_data    [0:`PE_COL-1][0:`W_C_LENGTH-1]; 
            logic        [`W_C_BITWIDTH-1:0]       i_w_c_idx   [0:`PE_COL-1][0:`W_C_LENGTH-1];
            logic        [`W_POS_PTR_BITWIDTH-1:0] i_pos_ptr   [0:`PE_COL-1][0:`W_R_LENGTH-1];
            logic        [`W_R_BITWIDTH-1:0]       i_r_idx     [0:`PE_COL-1][0:`W_R_LENGTH-1];
            logic        [`W_K_BITWIDTH-1:0]       i_k_idx     [0:`PE_COL-1][0:`W_R_LENGTH-1];
            logic        [1:0]                     i_w_s       [0:`PE_COL-1];
            logic        [$clog2(`W_C_LENGTH):0] i_w_iters   [0:`PE_COL-1];
            logic        [$clog2(`W_C_LENGTH):0] i_w_len     [0:`PE_COL-1];

            // Output
            logic                                  o_finish_PE [0:`PE_ROW-1][0:`PE_COL-1];
            logic signed [`IA_DATA_BITWIDTH-1:0]   o_OA        [0:`PE_ROW-1][0:`PE_COL-1][0:`IA_ROW*`IA_CHANNEL-1];
            
        // ----------------------- Else ------------------------
            logic                                  o_finish_CAMERA;
            

    // ========================== Logic (Reg) =============================
        // For PE
        logic                                   i_start_PEs, i_start_PEs_n;
        logic        [$clog2(`IA_CHANNEL):0]  ia_iters    [0:`IA_ROW-1][0:`IA_COL-1],                  ia_iters_n    [0:`IA_ROW-1][0:`IA_COL-1];
        logic        [$clog2(`IA_CHANNEL):0]  ia_len      [0:`IA_ROW-1][0:`IA_COL-1],                  ia_len_n      [0:`IA_ROW-1][0:`IA_COL-1];
        // For OA
        logic signed [`IA_DATA_BITWIDTH-1:0]    oa_buffer   [0:`IA_ROW-1][0:`IA_COL-1][0:`IA_CHANNEL-1], oa_buffer_n   [0:`IA_ROW-1][0:`IA_COL-1][0:`IA_CHANNEL-1];
        logic signed [`IA_DATA_BITWIDTH-1:0]    oa_reducer  [0:`IA_ROW+`IA_COL-2][0:2][0:`IA_CHANNEL-1], oa_reducer_n  [0:`IA_ROW+`IA_COL-2][0:2][0:`IA_CHANNEL-1];
        logic signed [`IA_DATA_BITWIDTH-1:0]    ia_data     [0:`IA_ROW-1][0:`IA_COL-1][0:`IA_CHANNEL-1], ia_data_n     [0:`IA_ROW-1][0:`IA_COL-1][0:`IA_CHANNEL-1];
        logic        [`IA_C_BITWIDTH-1:0]       ia_c_idx    [0:`IA_ROW-1][0:`IA_COL-1][0:`IA_CHANNEL-1], ia_c_idx_n    [0:`IA_ROW-1][0:`IA_COL-1][0:`IA_CHANNEL-1];
        logic        [4:0]                      state, state_n;
        logic        [$clog2(`IA_ROW) :0]      Hi, Hi_n,                  h, h_n;
        logic        [$clog2(`IA_COL) :0]      Wi, Wi_n,                  w_start_max, w_start_max_n,      w_start, w_start_n;        
        logic        [$clog2(`IA_CHANNEL):0]  Co, Co_n;

        // Maxpool


    // ========================== PE Arrays (7 x 3) === unfinished ==========================
        generate
            for (genvar gv_row=0; gv_row < `PE_ROW; gv_row++) begin
                for (genvar gv_col=0; gv_col < `PE_COL; gv_col++) begin
                    PE_TEMP u_PE_TEMP(
                        .i_clk          (i_clk),
                        .i_rst_n        (i_rst_n),
                        .i_start        (i_start_PEs),
                        // IA bundle
                        .i_ia_h         (i_ia_h    [gv_row]),
                        .i_ia_w         (i_ia_w    [gv_row]),
                        .i_ia_data      (i_ia_data [gv_row]),
                        .i_ia_c_idx     (i_ia_c_idx[gv_row]),
                        .i_ia_iters     (i_ia_iters[gv_row]),
                        .i_ia_len       (i_ia_len  [gv_row]),
                        // W bundle
                        .i_w_s          (i_w_s      [gv_col]),
                        .i_w_data       (i_w_data   [gv_col]),
                        .i_w_c_idx      (i_w_c_idx  [gv_col]),
                        .i_pos_ptr      (i_pos_ptr  [gv_col]),
                        .i_r_idx        (i_r_idx    [gv_col]),
                        .i_k_idx        (i_k_idx    [gv_col]),
                        .i_w_iters      (i_w_iters  [gv_col]),
                        .i_w_len        (i_w_len    [gv_col]),

                        // Output
                        .o_finish       (o_finish_PE[gv_row][gv_col]),
                        .o_OA           (o_OA[gv_row][gv_col])
                    );
                end
            end
        endgenerate


    // ========================== Task ==================================================
        // task READ_i_w_data;
            
        // endtask
        task PUT_W;
            // remenber to reset all buffer except IA
            for (int r=0; r < `IA_ROW; r++ ) begin
                for (int c=0; c < `IA_COL; c++ ) begin
                    for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                        oa_buffer_n[r][c][ch] = 0;
                    end
                end
            end

            for (int id=0; id < `IA_ROW+`IA_COL-2; id++ ) begin
                for (int row=0; row < 3; row++ ) begin
                    for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                        oa_reducer_n[id][row][ch] = 0;
                    end
                end
            end

            case(state)
                S_PUT_W_1: begin

                    // 
                    for (int k=0; k < `W_C_LENGTH; k++) begin
                            i_w_data[0][k]    = (k<`W_C_LENGTH_L1_S0) ? $signed( w_data_l1_s0[k] ) : -1;
                            i_w_data[1][k]    = (k<`W_C_LENGTH_L1_S1) ? $signed( w_data_l1_s1[k] ) : -1;
                            i_w_data[2][k]    = (k<`W_C_LENGTH_L1_S2) ? $signed( w_data_l1_s2[k] ) : -1;

                            i_w_c_idx[0][k]   = (k<`W_C_LENGTH_L1_S0) ?          w_c_idx_l1_s0[k]   : 0; 
                            i_w_c_idx[1][k]   = (k<`W_C_LENGTH_L1_S1) ?          w_c_idx_l1_s1[k]   : 0; 
                            i_w_c_idx[2][k]   = (k<`W_C_LENGTH_L1_S2) ?          w_c_idx_l1_s2[k]   : 0; 

                            i_pos_ptr[0][k]   = (k<`W_R_LENGTH_L1_S0) ?          w_pos_ptr_l1_s0[k] : 0; 
                            i_pos_ptr[1][k]   = (k<`W_R_LENGTH_L1_S1) ?          w_pos_ptr_l1_s1[k] : 0; 
                            i_pos_ptr[2][k]   = (k<`W_R_LENGTH_L1_S2) ?          w_pos_ptr_l1_s2[k] : 0; 


                            i_r_idx[0][k]     = (k<`W_R_LENGTH_L1_S0) ?          w_r_idx_l1_s0[k]   : 0; 
                            i_r_idx[1][k]     = (k<`W_R_LENGTH_L1_S1) ?          w_r_idx_l1_s1[k]   : 0; 
                            i_r_idx[2][k]     = (k<`W_R_LENGTH_L1_S2) ?          w_r_idx_l1_s2[k]   : 0; 

                            i_k_idx[0][k]     = (k<`W_R_LENGTH_L1_S0) ?          w_k_idx_l1_s0[k]   : 0; 
                            i_k_idx[1][k]     = (k<`W_R_LENGTH_L1_S1) ?          w_k_idx_l1_s1[k]   : 0; 
                            i_k_idx[2][k]     = (k<`W_R_LENGTH_L1_S2) ?          w_k_idx_l1_s2[k]   : 0; 
                    end
            

                    for (int pe_col=0; pe_col < `PE_COL; pe_col++) begin 
                        i_w_s       [pe_col] = w_s          [pe_col];
                        i_w_len     [pe_col] = w_len_1      [pe_col];
                        i_w_iters   [pe_col] = w_iters_1    [pe_col];
                    end

                    



                end

                S_PUT_W_2: begin
                    // 
                    for (int k=0; k < `W_C_LENGTH; k++) begin
                            i_w_data[0][k]    = (k<`W_C_LENGTH_L2_S0) ? $signed( w_data_l2_s0[k] ) : -1;
                            i_w_data[1][k]    = (k<`W_C_LENGTH_L2_S1) ? $signed( w_data_l2_s1[k] ) : -1;
                            i_w_data[2][k]    = (k<`W_C_LENGTH_L2_S2) ? $signed( w_data_l2_s2[k] ) : -1;

                            i_w_c_idx[0][k]   = (k<`W_C_LENGTH_L2_S0) ?          w_c_idx_l2_s0[k]   : 0; 
                            i_w_c_idx[1][k]   = (k<`W_C_LENGTH_L2_S1) ?          w_c_idx_l2_s1[k]   : 0; 
                            i_w_c_idx[2][k]   = (k<`W_C_LENGTH_L2_S2) ?          w_c_idx_l2_s2[k]   : 0; 

                            i_pos_ptr[0][k]   = (k<`W_R_LENGTH_L2_S0) ?          w_pos_ptr_l2_s0[k] : 0; 
                            i_pos_ptr[1][k]   = (k<`W_R_LENGTH_L2_S1) ?          w_pos_ptr_l2_s1[k] : 0; 
                            i_pos_ptr[2][k]   = (k<`W_R_LENGTH_L2_S2) ?          w_pos_ptr_l2_s2[k] : 0; 


                            i_r_idx[0][k]     = (k<`W_R_LENGTH_L2_S0) ?          w_r_idx_l2_s0[k]   : 0; 
                            i_r_idx[1][k]     = (k<`W_R_LENGTH_L2_S1) ?          w_r_idx_l2_s1[k]   : 0; 
                            i_r_idx[2][k]     = (k<`W_R_LENGTH_L2_S2) ?          w_r_idx_l2_s2[k]   : 0; 

                            i_k_idx[0][k]     = (k<`W_R_LENGTH_L2_S0) ?          w_k_idx_l2_s0[k]   : 0; 
                            i_k_idx[1][k]     = (k<`W_R_LENGTH_L2_S1) ?          w_k_idx_l2_s1[k]   : 0; 
                            i_k_idx[2][k]     = (k<`W_R_LENGTH_L2_S2) ?          w_k_idx_l2_s2[k]   : 0; 
                    end
            
                    for (int pe_col=0; pe_col < `PE_COL; pe_col++) begin 
                        i_w_s       [pe_col] = w_s          [pe_col];
                        i_w_len     [pe_col] = w_len_2      [pe_col];
                        i_w_iters   [pe_col] = w_iters_2    [pe_col];
                    end

                    
                    
                end
            endcase
        endtask


        task CONV;    // finish
            i_start_PEs_n = 1;
            for (int pe_row=0; pe_row < `PE_ROW; pe_row++) begin 
                i_ia_h      [pe_row]  =         h;
                i_ia_w      [pe_row]  =         w_start + pe_row;
                i_ia_data   [pe_row]  = $signed(ia_data     [h][w_start + pe_row] );
                i_ia_c_idx  [pe_row]  =         ia_c_idx    [h][w_start + pe_row];
                i_ia_iters  [pe_row]  =         ia_iters    [h][w_start + pe_row];
                i_ia_len    [pe_row]  =         ia_len      [h][w_start + pe_row];
            end
        endtask

        task TOOABUFFER;   
            // didn;t write code like : " (ch < Co ) ? ... :... ", Since I think  it need not to do,  Just to handle Co  when Compression or next layer's Hi

            // input [$clog2(`IA_COL)-1:0] w_start;
            // input [$clog2(`IA_ROW)-1:0] h;
            case(w_start)
                0:  begin
                    case(h)
                        0: begin
                            for (int c=0; c < `PE_ROW; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[0][c][ch] = $signed(oa_buffer[0][c][ch]) + $signed(oa_reducer[c+2][2][ch]);
                                end
                            end
                        end
                        1: begin
                            for (int c=0; c < `PE_ROW; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[0][c][ch] = $signed(oa_buffer[0][c][ch]) + $signed(oa_reducer[c+2][1][ch]);
                                    oa_buffer_n[1][c][ch] = $signed(oa_buffer[1][c][ch]) + $signed(oa_reducer[c+2][2][ch]);
                                end
                            end    
                        end
                        (Hi-2): begin
                            for (int c=0; c < `PE_ROW; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c+2][0][ch]);
                                    oa_buffer_n[h-1][c][ch] = $signed(oa_buffer[h-1][c][ch]) + $signed(oa_reducer[c+2][1][ch]);
                                end
                            end                              
                        end
                        (Hi-1): begin
                            for (int c=0; c < `PE_ROW; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c+2][0][ch]);
                                end
                            end 
                        end
                        default: begin
                            for (int c=0; c < `PE_ROW; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c+2][0][ch]);
                                    oa_buffer_n[h-1][c][ch] = $signed(oa_buffer[h-1][c][ch]) + $signed(oa_reducer[c+2][1][ch]);
                                    oa_buffer_n[h  ][c][ch] = $signed(oa_buffer[h  ][c][ch]) + $signed(oa_reducer[c+2][2][ch]);
                                end
                            end  
                        end
                    endcase
                end
                (w_start_max-1):    begin
                    case(h)
                        0: begin
                            for (int c=w_start*7-2; c < Wi-1; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[0][c][ch] = $signed(oa_buffer[0][c][ch]) + $signed(oa_reducer[c-w_start*7+2][2][ch]);
                                end
                            end
                        end
                        1: begin
                            for (int c=w_start*7-2; c < Wi-1; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[0][c][ch] = $signed(oa_buffer[0][c][ch]) + $signed(oa_reducer[c-w_start*7+2][1][ch]);
                                    oa_buffer_n[1][c][ch] = $signed(oa_buffer[1][c][ch]) + $signed(oa_reducer[c-w_start*7+2][2][ch]);
                                end
                            end    
                        end
                        (Hi-2): begin
                            for (int c=w_start*7-2; c < Wi-1; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c-w_start*7+2][0][ch]);
                                    oa_buffer_n[h-1][c][ch] = $signed(oa_buffer[h-1][c][ch]) + $signed(oa_reducer[c-w_start*7+2][1][ch]);
                                end
                            end                              
                        end
                        (Hi-1): begin
                            for (int c=w_start*7-2; c < Wi-1; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c-w_start*7+2][0][ch]);
                                end
                            end 
                        end
                        default: begin
                            for (int c=w_start*7-2; c < Wi-1; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c-w_start*7+2][0][ch]);
                                    oa_buffer_n[h-1][c][ch] = $signed(oa_buffer[h-1][c][ch]) + $signed(oa_reducer[c-w_start*7+2][1][ch]);
                                    oa_buffer_n[h  ][c][ch] = $signed(oa_buffer[h  ][c][ch]) + $signed(oa_reducer[c-w_start*7+2][2][ch]);
                                end
                            end  
                        end
                    endcase
                end
                default:    begin
                     case(h)
                        0: begin
                            for (int c=w_start*7-2; c < w_start*7+7; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[0][c][ch] = $signed(oa_buffer[0][c][ch]) + $signed(oa_reducer[c-w_start*7+2][2][ch]);
                                end
                            end
                        end
                        1: begin
                            for (int c=w_start*7-2; c < w_start*7+7; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[0][c][ch] = $signed(oa_buffer[0][c][ch]) + $signed(oa_reducer[c-w_start*7+2][1][ch]);
                                    oa_buffer_n[1][c][ch] = $signed(oa_buffer[1][c][ch]) + $signed(oa_reducer[c-w_start*7+2][2][ch]);
                                end
                            end    
                        end
                        (Hi-2): begin
                            for (int c=w_start*7-2; c < w_start*7+7; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c-w_start*7+2][0][ch]);
                                    oa_buffer_n[h-1][c][ch] = $signed(oa_buffer[h-1][c][ch]) + $signed(oa_reducer[c-w_start*7+2][1][ch]);
                                end
                            end                              
                        end
                        (Hi-1): begin
                            for (int c=w_start*7-2; c < w_start*7+7; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c-w_start*7+2][0][ch]);
                                end
                            end 
                        end
                        default: begin
                            for (int c=w_start*7-2; c < w_start*7+7; c++ ) begin
                                for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                                    oa_buffer_n[h-2][c][ch] = $signed(oa_buffer[h-2][c][ch]) + $signed(oa_reducer[c-w_start*7+2][0][ch]);
                                    oa_buffer_n[h-1][c][ch] = $signed(oa_buffer[h-1][c][ch]) + $signed(oa_reducer[c-w_start*7+2][1][ch]);
                                    oa_buffer_n[h  ][c][ch] = $signed(oa_buffer[h  ][c][ch]) + $signed(oa_reducer[c-w_start*7+2][2][ch]);
                                end
                            end  
                        end
                    endcase
                end
            endcase
        endtask

        task TOOAREDUCER; // todo
            // Co
            for(int r=0; r<3; r++) begin
                for(int ch = 0; ch < `IA_CHANNEL; ch++) begin
                    oa_reducer_n[0][r][ch] = (ch < Co) ? $signed(o_OA[0][2][ Co*(2-r)+ch ])                                        : 0;
                    oa_reducer_n[1][r][ch] = (ch < Co) ? $signed(o_OA[0][1][ Co*(2-r)+ch ]) +  $signed(o_OA[1][2][ Co*(2-r)+ch ])  : 0;
                    oa_reducer_n[7][r][ch] = (ch < Co) ? $signed(o_OA[5][0][ Co*(2-r)+ch ]) +  $signed(o_OA[6][1][ Co*(2-r)+ch ])  : 0;
                    oa_reducer_n[8][r][ch] = (ch < Co) ? $signed(o_OA[6][0][ Co*(2-r)+ch ])                                        : 0;
                end
            end

            for (int id=2; id<7; id++ ) begin
                for(int r=0; r<3; r++) begin
                    for(int ch = 0; ch < `IA_CHANNEL; ch++) begin
                        oa_reducer_n[id][r][ch] = (ch < Co) ? $signed(o_OA[id-2][0][ Co*(2-r)+ch ]) +  $signed(o_OA[id-1][1][ Co*(2-r)+ch ]) +  $signed(o_OA[id][2][ Co*(2-r)+ch ])  : 0;                
                    end
                end
            end
        endtask 

        task COMPRESS;

        endtask

        task MAXPOOL;
            // for (int r=0; r< (`IA))

        endtask

    // ========================== State Control (Combinational Circuit) ========= unfinish============
        always_comb begin  
            state_n = state;
            case(state)
                S_IDLE:         state_n = (i_start)                   ? S_CAMERA : state;
                // S_CAMERA:       state_n = (o_finish_CAMERA)           ? S_PUT_W_1 : state;
                // S_IDLE:         state_n = S_CAMERA;
                S_CAMERA:       state_n = S_PUT_W_1;
                S_PUT_W_1:      state_n = S_CONV_1;
                S_CONV_1:       state_n = (o_finish_PE==PEs_FINISH)   ? S_REDUCE_1 : state; 
                S_REDUCE_1:     state_n = S_TOOABUFFER_1;
                S_TOOABUFFER_1: state_n = (h==Hi-1 && w_start==w_start_max-1) ? S_COMPRESS_1 : S_CONV_1;

                S_COMPRESS_1:   state_n = S_PUT_W_2; // need to rethink

                S_PUT_W_2:      state_n = S_CONV_2;
                S_CONV_2:       state_n = (o_finish_PE==PEs_FINISH)   ? S_REDUCE_2 : state; 
                S_REDUCE_2:     state_n = S_TOOABUFFER_2;
                S_TOOABUFFER_2:       state_n = (h==Hi-1 && w_start==w_start_max-1) ? S_MAXPOOL  : S_CONV_2;

                S_MAXPOOL:      state_n = S_LINEAR; // need to rethink
                S_LINEAR:       state_n = S_OUT;    // need to rethink
                // S_OUT:          state_n = S_CAMERA; // need to rethink

                
            endcase
        end


    // ========================== Combinational Circuit =====unfinish================================
        always_comb begin 
            i_start_PEs_n  = i_start_PEs;
            o_random_out_n = o_random_out;
            Hi_n           = Hi;
            Wi_n           = Wi;
            w_start_max_n  = w_start_max;
            h_n            = h;
            w_start_n      = w_start;
            Co_n           = Co;

            ia_iters_n     = ia_iters;
            ia_len_n       = ia_len;
            ia_data_n      = ia_data;
            ia_c_idx_n     = ia_c_idx;
            oa_reducer_n   = oa_reducer;
            oa_buffer_n    = oa_buffer;

            case(state)
                S_IDLE: begin
                end

                S_CAMERA: begin
                end

                S_PUT_W_1: begin
                    PUT_W();
                    Hi_n = 16;
                    Wi_n = 16;
                    Co_n = 8;
                    w_start_max_n = 3;
                end

                S_CONV_1 : begin
                    CONV();

                end

                S_REDUCE_1: begin
                    TOOAREDUCER();
                    i_start_PEs_n = 0;
                end

                S_TOOABUFFER_1: begin // put to oa_buffer
                    TOOABUFFER();
                    h_n = (h == Hi-1) ? 0 : h+1;
                    if (h==Hi-1) begin
                        w_start_n = (w_start == w_start_max-1) ? 0 : w_start+1;
                    end
                end

                S_COMPRESS_1: begin // put to IA
                end

                S_PUT_W_2: begin
                    PUT_W();
                    Hi_n = 14;
                    Wi_n = 14;
                    Co_n = 8;
                    w_start_max_n = 2;
                end

                S_CONV_2 : begin
                    CONV();
                end

                S_REDUCE_2: begin
                    TOOAREDUCER();
                    i_start_PEs_n = 0;
                end

                S_TOOABUFFER_2: begin // put to oa_buffer
                    TOOABUFFER();
                    h_n = (h == Hi-1) ? 0 : h+1;
                    if (h==Hi-1) begin
                        w_start_n = (w_start == w_start_max-1) ? 0 : w_start+1;
                    end
                end

                S_MAXPOOL: begin // from oa_buffer to ia_buffer, one cycle
                end

                S_LINEAR : begin
                end

                S_OUT    : begin
                end

            endcase

        end

    // ========================== Sequential Circuit ========================================
        always_ff @(posedge i_clk or negedge i_rst_n) begin
            if (!i_rst_n) begin
                i_start_PEs  <= 0;
                o_random_out <= 0;
                state        <= S_IDLE;
                Hi           <= 0;
                Wi           <= 0;
                w_start_max  <= 0;
                h            <= 0;
                w_start      <= 0;
                Co           <= 0;

                

                for (int r=0; r < `IA_ROW; r++ ) begin
                    for (int c=0; c < `IA_COL; c++ ) begin
                        ia_iters [r][c] <= 0;
                        ia_len   [r][c] <= 0;
                        for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                            ia_data  [r][c][ch] <= 0;
                            ia_c_idx [r][c][ch] <= 0;
                            oa_buffer[r][c][ch] <= 0;
                        end
                    end
                end

                for (int id=0; id < `IA_ROW+`IA_COL-2; id++ ) begin
                    for (int row=0; row < 3; row++ ) begin
                        for (int ch=0; ch < `IA_CHANNEL; ch++ ) begin
                            oa_reducer[id][row][ch] <= 0;
                        end
                    end
                end

                
            end
            else begin
                i_start_PEs  <= i_start_PEs_n;
                o_random_out <= o_random_out_n;
                state        <= state_n;
                Hi           <= Hi_n;
                Wi           <= Wi_n;
                w_start_max  <= w_start_max_n;
                h            <= h_n;
                w_start      <= w_start_n;
                Co           <= Co_n;

                ia_iters     <= ia_iters_n;
                ia_len       <= ia_len_n;
                ia_data      <= ia_data_n;
                ia_c_idx     <= ia_c_idx_n;
                oa_reducer   <= oa_reducer_n;
                oa_buffer    <= oa_buffer_n;
                

            end

        end

endmodule

















