// w_data
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_DATA_BITWIDTH'b1111110011100101,
        `W_DATA_BITWIDTH'b1111111001011110,
        `W_DATA_BITWIDTH'b0000001001011101,
        `W_DATA_BITWIDTH'b1111111101011000,
        `W_DATA_BITWIDTH'b1111110101101101,
        `W_DATA_BITWIDTH'b1111110010110110,
        `W_DATA_BITWIDTH'b0000001110111010,
        `W_DATA_BITWIDTH'b1111111010001100,
        `W_DATA_BITWIDTH'b0000001000001011,
        `W_DATA_BITWIDTH'b1111101111110111,
        `W_DATA_BITWIDTH'b0000000010111010,
        `W_DATA_BITWIDTH'b0000001101011100,
        `W_DATA_BITWIDTH'b0000000110001011,
        `W_DATA_BITWIDTH'b1111110000101100,
        `W_DATA_BITWIDTH'b0000001110000100,
        `W_DATA_BITWIDTH'b0000010011010001,
        `W_DATA_BITWIDTH'b1111100001100110,
        `W_DATA_BITWIDTH'b0000001110000111,
        `W_DATA_BITWIDTH'b1111110110101001,
        `W_DATA_BITWIDTH'b1111111000011000,
        `W_DATA_BITWIDTH'b0000001000010001,
        `W_DATA_BITWIDTH'b0000000110110111,
        `W_DATA_BITWIDTH'b0000000010000000,
        `W_DATA_BITWIDTH'b1111110100000000,
        `W_DATA_BITWIDTH'b0000000110010101,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b0000000101011011,
        `W_DATA_BITWIDTH'b0000001000101100,
        `W_DATA_BITWIDTH'b0000000111010100,
        `W_DATA_BITWIDTH'b1111111000001000,
        `W_DATA_BITWIDTH'b1111111011011010,
        `W_DATA_BITWIDTH'b0000000010011110,
        `W_DATA_BITWIDTH'b1111111100110001,
        `W_DATA_BITWIDTH'b0000010000101111,
        `W_DATA_BITWIDTH'b1111101001000011,
        `W_DATA_BITWIDTH'b1111111000011101,
        `W_DATA_BITWIDTH'b1111110010111111,
        `W_DATA_BITWIDTH'b1111111101110010,
        `W_DATA_BITWIDTH'b1111111011110001,
        `W_DATA_BITWIDTH'b1111111011100011,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000111100110,
        `W_DATA_BITWIDTH'b0000010001100000,
        `W_DATA_BITWIDTH'b1111101101100010,
        `W_DATA_BITWIDTH'b1111111101110110,
        `W_DATA_BITWIDTH'b0000001110000101,
        `W_DATA_BITWIDTH'b1111100111001110,
        `W_DATA_BITWIDTH'b0000000101011000,
        `W_DATA_BITWIDTH'b0000001101011101,
        `W_DATA_BITWIDTH'b1111110000000010,
        `W_DATA_BITWIDTH'b0000001000001000,
        `W_DATA_BITWIDTH'b1111100111110100,
        `W_DATA_BITWIDTH'b0000000111100011,
        `W_DATA_BITWIDTH'b0000001001010101,
        `W_DATA_BITWIDTH'b0000000100011010,
        `W_DATA_BITWIDTH'b0000010011000111,
        `W_DATA_BITWIDTH'b0000000010000001,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000000011100001,
        `W_DATA_BITWIDTH'b1111111010100101,
        `W_DATA_BITWIDTH'b0000000101001001,
        `W_DATA_BITWIDTH'b0000001111100110,
        `W_DATA_BITWIDTH'b0000001010101001,
        `W_DATA_BITWIDTH'b0000011011010011,
        `W_DATA_BITWIDTH'b1111101100010100,
        `W_DATA_BITWIDTH'b0000000010010101,
        `W_DATA_BITWIDTH'b1111101001100110,
        `W_DATA_BITWIDTH'b1111101001100110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_DATA_BITWIDTH'b0000001011111110,
        `W_DATA_BITWIDTH'b0000000001111100,
        `W_DATA_BITWIDTH'b0000000100001101,
        `W_DATA_BITWIDTH'b0000001001111011,
        `W_DATA_BITWIDTH'b1111111011100110,
        `W_DATA_BITWIDTH'b1111111010000111,
        `W_DATA_BITWIDTH'b1111101111000001,
        `W_DATA_BITWIDTH'b1111111101100001,
        `W_DATA_BITWIDTH'b0000011011100110,
        `W_DATA_BITWIDTH'b0000000011100101,
        `W_DATA_BITWIDTH'b1111110011101111,
        `W_DATA_BITWIDTH'b0000000011101000,
        `W_DATA_BITWIDTH'b1111110100010101,
        `W_DATA_BITWIDTH'b1111110010010100,
        `W_DATA_BITWIDTH'b1111110011100001,
        `W_DATA_BITWIDTH'b0000000101010100,
        `W_DATA_BITWIDTH'b1111110111011100,
        `W_DATA_BITWIDTH'b1111110111011000,
        `W_DATA_BITWIDTH'b0000000101001100,
        `W_DATA_BITWIDTH'b1111110100010011,
        `W_DATA_BITWIDTH'b1111111010011111,
        `W_DATA_BITWIDTH'b0000001001100101,
        `W_DATA_BITWIDTH'b0000000111010101,
        `W_DATA_BITWIDTH'b1111100101110011,
        `W_DATA_BITWIDTH'b0000011010010111,
        `W_DATA_BITWIDTH'b0000000011000011,
        `W_DATA_BITWIDTH'b1111110101101010,
        `W_DATA_BITWIDTH'b0000000110111011,
        `W_DATA_BITWIDTH'b1111101110111011,
        `W_DATA_BITWIDTH'b0000010111100100,
        `W_DATA_BITWIDTH'b0000000110001111,
        `W_DATA_BITWIDTH'b0000010000001011,
        `W_DATA_BITWIDTH'b1111110111001100,
        `W_DATA_BITWIDTH'b1111111001100010,
        `W_DATA_BITWIDTH'b0000000101110101,
        `W_DATA_BITWIDTH'b1111101101101110,
        `W_DATA_BITWIDTH'b0000000100001110,
        `W_DATA_BITWIDTH'b0000000110111001,
        `W_DATA_BITWIDTH'b1111111100110110,
        `W_DATA_BITWIDTH'b1111111100101010,
        `W_DATA_BITWIDTH'b0000000111111111,
        `W_DATA_BITWIDTH'b0000100101101101,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110000000101,
        `W_DATA_BITWIDTH'b1111110000011011,
        `W_DATA_BITWIDTH'b0000000010110101,
        `W_DATA_BITWIDTH'b0000011010110011,
        `W_DATA_BITWIDTH'b1111111001101110,
        `W_DATA_BITWIDTH'b0000000101011110,
        `W_DATA_BITWIDTH'b1111111011001011,
        `W_DATA_BITWIDTH'b0000001101111000,
        `W_DATA_BITWIDTH'b0000011010000001,
        `W_DATA_BITWIDTH'b1111100010110110,
        `W_DATA_BITWIDTH'b1111110111010110,
        `W_DATA_BITWIDTH'b0000011010111110,
        `W_DATA_BITWIDTH'b1111101110100010,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b0000001000000110,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111100010100101,
        `W_DATA_BITWIDTH'b1111111011100000,
        `W_DATA_BITWIDTH'b0000001110100010,
        `W_DATA_BITWIDTH'b0000000111011111,
        `W_DATA_BITWIDTH'b1111110010111011,
        `W_DATA_BITWIDTH'b0000010000100101,
        `W_DATA_BITWIDTH'b0000010000100101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_DATA_BITWIDTH'b1111111101010101,
        `W_DATA_BITWIDTH'b0000000011101111,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110101011010,
        `W_DATA_BITWIDTH'b1111110101010100,
        `W_DATA_BITWIDTH'b0000001011110011,
        `W_DATA_BITWIDTH'b1111111001100101,
        `W_DATA_BITWIDTH'b0000010101111110,
        `W_DATA_BITWIDTH'b0000010010100101,
        `W_DATA_BITWIDTH'b1111011110010000,
        `W_DATA_BITWIDTH'b1111110001000001,
        `W_DATA_BITWIDTH'b0000001101001011,
        `W_DATA_BITWIDTH'b0000011001011010,
        `W_DATA_BITWIDTH'b1111100001111110,
        `W_DATA_BITWIDTH'b0000010010100111,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b1111111000111101,
        `W_DATA_BITWIDTH'b1111111011111100,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000110001000,
        `W_DATA_BITWIDTH'b1111110011001010,
        `W_DATA_BITWIDTH'b1111111001000011,
        `W_DATA_BITWIDTH'b1111111001011001,
        `W_DATA_BITWIDTH'b0000001010000101,
        `W_DATA_BITWIDTH'b0000001100001100,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111111001001011,
        `W_DATA_BITWIDTH'b0000010001001101,
        `W_DATA_BITWIDTH'b0000100000011111,
        `W_DATA_BITWIDTH'b1111100000100000,
        `W_DATA_BITWIDTH'b1111100111110111,
        `W_DATA_BITWIDTH'b0000001011100001,
        `W_DATA_BITWIDTH'b1111111101101011,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b0000001010100100,
        `W_DATA_BITWIDTH'b1111111000111110,
        `W_DATA_BITWIDTH'b0000001000000011,
        `W_DATA_BITWIDTH'b1111110101011011,
        `W_DATA_BITWIDTH'b1111111011010100,
        `W_DATA_BITWIDTH'b0000010010110001,
        `W_DATA_BITWIDTH'b1111110110001010,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b0000001110100101,
        `W_DATA_BITWIDTH'b0000000011100100,
        `W_DATA_BITWIDTH'b0000000111101001,
        `W_DATA_BITWIDTH'b0000001110011000,
        `W_DATA_BITWIDTH'b1111111101101010,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000001100101010,
        `W_DATA_BITWIDTH'b0000001001011111,
        `W_DATA_BITWIDTH'b1111111001010011,
        `W_DATA_BITWIDTH'b1111101010010111,
        `W_DATA_BITWIDTH'b1111110010010011,
        `W_DATA_BITWIDTH'b0000001111110100,
        `W_DATA_BITWIDTH'b0000000111011011,
        `W_DATA_BITWIDTH'b0000001011110101,
        `W_DATA_BITWIDTH'b1111100111101101,
        `W_DATA_BITWIDTH'b0000100000011000,
        `W_DATA_BITWIDTH'b1111111011111101,
        `W_DATA_BITWIDTH'b1111111011111101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_DATA_BITWIDTH'b1111110011100101,
        `W_DATA_BITWIDTH'b1111111001011110,
        `W_DATA_BITWIDTH'b0000001001011101,
        `W_DATA_BITWIDTH'b1111111101011000,
        `W_DATA_BITWIDTH'b1111110101101101,
        `W_DATA_BITWIDTH'b1111110010110110,
        `W_DATA_BITWIDTH'b0000001110111010,
        `W_DATA_BITWIDTH'b1111111010001100,
        `W_DATA_BITWIDTH'b0000001000001011,
        `W_DATA_BITWIDTH'b1111101111110111,
        `W_DATA_BITWIDTH'b0000000010111010,
        `W_DATA_BITWIDTH'b0000001101011100,
        `W_DATA_BITWIDTH'b0000000110001011,
        `W_DATA_BITWIDTH'b1111110000101100,
        `W_DATA_BITWIDTH'b0000001110000100,
        `W_DATA_BITWIDTH'b0000010011010001,
        `W_DATA_BITWIDTH'b1111100001100110,
        `W_DATA_BITWIDTH'b0000001110000111,
        `W_DATA_BITWIDTH'b1111110110101001,
        `W_DATA_BITWIDTH'b1111111000011000,
        `W_DATA_BITWIDTH'b0000001000010001,
        `W_DATA_BITWIDTH'b0000000110110111,
        `W_DATA_BITWIDTH'b0000000010000000,
        `W_DATA_BITWIDTH'b1111110100000000,
        `W_DATA_BITWIDTH'b0000000110010101,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b0000000101011011,
        `W_DATA_BITWIDTH'b0000001000101100,
        `W_DATA_BITWIDTH'b0000000111010100,
        `W_DATA_BITWIDTH'b1111111000001000,
        `W_DATA_BITWIDTH'b1111111011011010,
        `W_DATA_BITWIDTH'b0000000010011110,
        `W_DATA_BITWIDTH'b1111111100110001,
        `W_DATA_BITWIDTH'b0000010000101111,
        `W_DATA_BITWIDTH'b1111101001000011,
        `W_DATA_BITWIDTH'b1111111000011101,
        `W_DATA_BITWIDTH'b1111110010111111,
        `W_DATA_BITWIDTH'b1111111101110010,
        `W_DATA_BITWIDTH'b1111111011110001,
        `W_DATA_BITWIDTH'b1111111011100011,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000111100110,
        `W_DATA_BITWIDTH'b0000010001100000,
        `W_DATA_BITWIDTH'b1111101101100010,
        `W_DATA_BITWIDTH'b1111111101110110,
        `W_DATA_BITWIDTH'b0000001110000101,
        `W_DATA_BITWIDTH'b1111100111001110,
        `W_DATA_BITWIDTH'b0000000101011000,
        `W_DATA_BITWIDTH'b0000001101011101,
        `W_DATA_BITWIDTH'b1111110000000010,
        `W_DATA_BITWIDTH'b0000001000001000,
        `W_DATA_BITWIDTH'b1111100111110100,
        `W_DATA_BITWIDTH'b0000000111100011,
        `W_DATA_BITWIDTH'b0000001001010101,
        `W_DATA_BITWIDTH'b0000000100011010,
        `W_DATA_BITWIDTH'b0000010011000111,
        `W_DATA_BITWIDTH'b0000000010000001,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000000011100001,
        `W_DATA_BITWIDTH'b1111111010100101,
        `W_DATA_BITWIDTH'b0000000101001001,
        `W_DATA_BITWIDTH'b0000001111100110,
        `W_DATA_BITWIDTH'b0000001010101001,
        `W_DATA_BITWIDTH'b0000011011010011,
        `W_DATA_BITWIDTH'b1111101100010100,
        `W_DATA_BITWIDTH'b0000000010010101,
        `W_DATA_BITWIDTH'b1111101001100110,
        `W_DATA_BITWIDTH'b1111101001100110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_DATA_BITWIDTH'b0000001011111110,
        `W_DATA_BITWIDTH'b0000000001111100,
        `W_DATA_BITWIDTH'b0000000100001101,
        `W_DATA_BITWIDTH'b0000001001111011,
        `W_DATA_BITWIDTH'b1111111011100110,
        `W_DATA_BITWIDTH'b1111111010000111,
        `W_DATA_BITWIDTH'b1111101111000001,
        `W_DATA_BITWIDTH'b1111111101100001,
        `W_DATA_BITWIDTH'b0000011011100110,
        `W_DATA_BITWIDTH'b0000000011100101,
        `W_DATA_BITWIDTH'b1111110011101111,
        `W_DATA_BITWIDTH'b0000000011101000,
        `W_DATA_BITWIDTH'b1111110100010101,
        `W_DATA_BITWIDTH'b1111110010010100,
        `W_DATA_BITWIDTH'b1111110011100001,
        `W_DATA_BITWIDTH'b0000000101010100,
        `W_DATA_BITWIDTH'b1111110111011100,
        `W_DATA_BITWIDTH'b1111110111011000,
        `W_DATA_BITWIDTH'b0000000101001100,
        `W_DATA_BITWIDTH'b1111110100010011,
        `W_DATA_BITWIDTH'b1111111010011111,
        `W_DATA_BITWIDTH'b0000001001100101,
        `W_DATA_BITWIDTH'b0000000111010101,
        `W_DATA_BITWIDTH'b1111100101110011,
        `W_DATA_BITWIDTH'b0000011010010111,
        `W_DATA_BITWIDTH'b0000000011000011,
        `W_DATA_BITWIDTH'b1111110101101010,
        `W_DATA_BITWIDTH'b0000000110111011,
        `W_DATA_BITWIDTH'b1111101110111011,
        `W_DATA_BITWIDTH'b0000010111100100,
        `W_DATA_BITWIDTH'b0000000110001111,
        `W_DATA_BITWIDTH'b0000010000001011,
        `W_DATA_BITWIDTH'b1111110111001100,
        `W_DATA_BITWIDTH'b1111111001100010,
        `W_DATA_BITWIDTH'b0000000101110101,
        `W_DATA_BITWIDTH'b1111101101101110,
        `W_DATA_BITWIDTH'b0000000100001110,
        `W_DATA_BITWIDTH'b0000000110111001,
        `W_DATA_BITWIDTH'b1111111100110110,
        `W_DATA_BITWIDTH'b1111111100101010,
        `W_DATA_BITWIDTH'b0000000111111111,
        `W_DATA_BITWIDTH'b0000100101101101,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110000000101,
        `W_DATA_BITWIDTH'b1111110000011011,
        `W_DATA_BITWIDTH'b0000000010110101,
        `W_DATA_BITWIDTH'b0000011010110011,
        `W_DATA_BITWIDTH'b1111111001101110,
        `W_DATA_BITWIDTH'b0000000101011110,
        `W_DATA_BITWIDTH'b1111111011001011,
        `W_DATA_BITWIDTH'b0000001101111000,
        `W_DATA_BITWIDTH'b0000011010000001,
        `W_DATA_BITWIDTH'b1111100010110110,
        `W_DATA_BITWIDTH'b1111110111010110,
        `W_DATA_BITWIDTH'b0000011010111110,
        `W_DATA_BITWIDTH'b1111101110100010,
        `W_DATA_BITWIDTH'b1111110101000100,
        `W_DATA_BITWIDTH'b0000001000000110,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111100010100101,
        `W_DATA_BITWIDTH'b1111111011100000,
        `W_DATA_BITWIDTH'b0000001110100010,
        `W_DATA_BITWIDTH'b0000000111011111,
        `W_DATA_BITWIDTH'b1111110010111011,
        `W_DATA_BITWIDTH'b0000010000100101,
        `W_DATA_BITWIDTH'b0000010000100101
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_DATA_BITWIDTH'b1111111101010101,
        `W_DATA_BITWIDTH'b0000000011101111,
        `W_DATA_BITWIDTH'b1111111100001011,
        `W_DATA_BITWIDTH'b1111110101011010,
        `W_DATA_BITWIDTH'b1111110101010100,
        `W_DATA_BITWIDTH'b0000001011110011,
        `W_DATA_BITWIDTH'b1111111001100101,
        `W_DATA_BITWIDTH'b0000010101111110,
        `W_DATA_BITWIDTH'b0000010010100101,
        `W_DATA_BITWIDTH'b1111011110010000,
        `W_DATA_BITWIDTH'b1111110001000001,
        `W_DATA_BITWIDTH'b0000001101001011,
        `W_DATA_BITWIDTH'b0000011001011010,
        `W_DATA_BITWIDTH'b1111100001111110,
        `W_DATA_BITWIDTH'b0000010010100111,
        `W_DATA_BITWIDTH'b1111110110111000,
        `W_DATA_BITWIDTH'b1111111000111101,
        `W_DATA_BITWIDTH'b1111111011111100,
        `W_DATA_BITWIDTH'b0000000110110011,
        `W_DATA_BITWIDTH'b0000000110001000,
        `W_DATA_BITWIDTH'b1111110011001010,
        `W_DATA_BITWIDTH'b1111111001000011,
        `W_DATA_BITWIDTH'b1111111001011001,
        `W_DATA_BITWIDTH'b0000001010000101,
        `W_DATA_BITWIDTH'b0000001100001100,
        `W_DATA_BITWIDTH'b1111111101100000,
        `W_DATA_BITWIDTH'b1111111001001011,
        `W_DATA_BITWIDTH'b0000010001001101,
        `W_DATA_BITWIDTH'b0000100000011111,
        `W_DATA_BITWIDTH'b1111100000100000,
        `W_DATA_BITWIDTH'b1111100111110111,
        `W_DATA_BITWIDTH'b0000001011100001,
        `W_DATA_BITWIDTH'b1111111101101011,
        `W_DATA_BITWIDTH'b1111111000111111,
        `W_DATA_BITWIDTH'b0000001010100100,
        `W_DATA_BITWIDTH'b1111111000111110,
        `W_DATA_BITWIDTH'b0000001000000011,
        `W_DATA_BITWIDTH'b1111110101011011,
        `W_DATA_BITWIDTH'b1111111011010100,
        `W_DATA_BITWIDTH'b0000010010110001,
        `W_DATA_BITWIDTH'b1111110110001010,
        `W_DATA_BITWIDTH'b1111110100001010,
        `W_DATA_BITWIDTH'b0000001110100101,
        `W_DATA_BITWIDTH'b0000000011100100,
        `W_DATA_BITWIDTH'b0000000111101001,
        `W_DATA_BITWIDTH'b0000001110011000,
        `W_DATA_BITWIDTH'b1111111101101010,
        `W_DATA_BITWIDTH'b1111101101100000,
        `W_DATA_BITWIDTH'b0000001100101010,
        `W_DATA_BITWIDTH'b0000001001011111,
        `W_DATA_BITWIDTH'b1111111001010011,
        `W_DATA_BITWIDTH'b1111101010010111,
        `W_DATA_BITWIDTH'b1111110010010011,
        `W_DATA_BITWIDTH'b0000001111110100,
        `W_DATA_BITWIDTH'b0000000111011011,
        `W_DATA_BITWIDTH'b0000001011110101,
        `W_DATA_BITWIDTH'b1111100111101101,
        `W_DATA_BITWIDTH'b0000100000011000,
        `W_DATA_BITWIDTH'b1111111011111101,
        `W_DATA_BITWIDTH'b1111111011111101
    };

// w_c_idx
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };
    localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00010,
        `W_C_BITWIDTH'b00000,
        `W_C_BITWIDTH'b00001,
        `W_C_BITWIDTH'b00001
    };

// w_r_idx
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };
    localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b10,
        `W_R_BITWIDTH'b00,
        `W_R_BITWIDTH'b01,
        `W_R_BITWIDTH'b01
    };

// w_k_idx
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };
    localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00000,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00001,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00010,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00011,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00100,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00101,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00110,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111,
        `W_K_BITWIDTH'b00111
    };

// w_pos_ptr
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000011,
        `W_POS_PTR_BITWIDTH'b00000000110,
        `W_POS_PTR_BITWIDTH'b00000001001,
        `W_POS_PTR_BITWIDTH'b00000001100,
        `W_POS_PTR_BITWIDTH'b00000001111,
        `W_POS_PTR_BITWIDTH'b00000010010,
        `W_POS_PTR_BITWIDTH'b00000010101,
        `W_POS_PTR_BITWIDTH'b00000011000,
        `W_POS_PTR_BITWIDTH'b00000011011,
        `W_POS_PTR_BITWIDTH'b00000011110,
        `W_POS_PTR_BITWIDTH'b00000100001,
        `W_POS_PTR_BITWIDTH'b00000100100,
        `W_POS_PTR_BITWIDTH'b00000100110,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000101010,
        `W_POS_PTR_BITWIDTH'b00000101101,
        `W_POS_PTR_BITWIDTH'b00000110000,
        `W_POS_PTR_BITWIDTH'b00000110011,
        `W_POS_PTR_BITWIDTH'b00000110110,
        `W_POS_PTR_BITWIDTH'b00000111001,
        `W_POS_PTR_BITWIDTH'b00000111011,
        `W_POS_PTR_BITWIDTH'b00000111110,
        `W_POS_PTR_BITWIDTH'b00000111110
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00001000100,
        `W_POS_PTR_BITWIDTH'b00001000111,
        `W_POS_PTR_BITWIDTH'b00001001001,
        `W_POS_PTR_BITWIDTH'b00001001100,
        `W_POS_PTR_BITWIDTH'b00001001111,
        `W_POS_PTR_BITWIDTH'b00001010001,
        `W_POS_PTR_BITWIDTH'b00001010100,
        `W_POS_PTR_BITWIDTH'b00001010111,
        `W_POS_PTR_BITWIDTH'b00001011000,
        `W_POS_PTR_BITWIDTH'b00001011011,
        `W_POS_PTR_BITWIDTH'b00001011110,
        `W_POS_PTR_BITWIDTH'b00001100001,
        `W_POS_PTR_BITWIDTH'b00001100100,
        `W_POS_PTR_BITWIDTH'b00001100111,
        `W_POS_PTR_BITWIDTH'b00001101010,
        `W_POS_PTR_BITWIDTH'b00001101101,
        `W_POS_PTR_BITWIDTH'b00001110000,
        `W_POS_PTR_BITWIDTH'b00001110011,
        `W_POS_PTR_BITWIDTH'b00001110110,
        `W_POS_PTR_BITWIDTH'b00001111001,
        `W_POS_PTR_BITWIDTH'b00001111100,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010000010,
        `W_POS_PTR_BITWIDTH'b00010000010
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00010000110,
        `W_POS_PTR_BITWIDTH'b00010001001,
        `W_POS_PTR_BITWIDTH'b00010001010,
        `W_POS_PTR_BITWIDTH'b00010001100,
        `W_POS_PTR_BITWIDTH'b00010001111,
        `W_POS_PTR_BITWIDTH'b00010010001,
        `W_POS_PTR_BITWIDTH'b00010010100,
        `W_POS_PTR_BITWIDTH'b00010010111,
        `W_POS_PTR_BITWIDTH'b00010011010,
        `W_POS_PTR_BITWIDTH'b00010011100,
        `W_POS_PTR_BITWIDTH'b00010011111,
        `W_POS_PTR_BITWIDTH'b00010100010,
        `W_POS_PTR_BITWIDTH'b00010100101,
        `W_POS_PTR_BITWIDTH'b00010100110,
        `W_POS_PTR_BITWIDTH'b00010101000,
        `W_POS_PTR_BITWIDTH'b00010101001,
        `W_POS_PTR_BITWIDTH'b00010101100,
        `W_POS_PTR_BITWIDTH'b00010101111,
        `W_POS_PTR_BITWIDTH'b00010110010,
        `W_POS_PTR_BITWIDTH'b00010110101,
        `W_POS_PTR_BITWIDTH'b00010110110,
        `W_POS_PTR_BITWIDTH'b00010111001,
        `W_POS_PTR_BITWIDTH'b00010111100,
        `W_POS_PTR_BITWIDTH'b00010111100
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000011,
        `W_POS_PTR_BITWIDTH'b00000000110,
        `W_POS_PTR_BITWIDTH'b00000001001,
        `W_POS_PTR_BITWIDTH'b00000001100,
        `W_POS_PTR_BITWIDTH'b00000001111,
        `W_POS_PTR_BITWIDTH'b00000010010,
        `W_POS_PTR_BITWIDTH'b00000010101,
        `W_POS_PTR_BITWIDTH'b00000011000,
        `W_POS_PTR_BITWIDTH'b00000011011,
        `W_POS_PTR_BITWIDTH'b00000011110,
        `W_POS_PTR_BITWIDTH'b00000100001,
        `W_POS_PTR_BITWIDTH'b00000100100,
        `W_POS_PTR_BITWIDTH'b00000100110,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000101010,
        `W_POS_PTR_BITWIDTH'b00000101101,
        `W_POS_PTR_BITWIDTH'b00000110000,
        `W_POS_PTR_BITWIDTH'b00000110011,
        `W_POS_PTR_BITWIDTH'b00000110110,
        `W_POS_PTR_BITWIDTH'b00000111001,
        `W_POS_PTR_BITWIDTH'b00000111011,
        `W_POS_PTR_BITWIDTH'b00000111110,
        `W_POS_PTR_BITWIDTH'b00000111110
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00001000100,
        `W_POS_PTR_BITWIDTH'b00001000111,
        `W_POS_PTR_BITWIDTH'b00001001001,
        `W_POS_PTR_BITWIDTH'b00001001100,
        `W_POS_PTR_BITWIDTH'b00001001111,
        `W_POS_PTR_BITWIDTH'b00001010001,
        `W_POS_PTR_BITWIDTH'b00001010100,
        `W_POS_PTR_BITWIDTH'b00001010111,
        `W_POS_PTR_BITWIDTH'b00001011000,
        `W_POS_PTR_BITWIDTH'b00001011011,
        `W_POS_PTR_BITWIDTH'b00001011110,
        `W_POS_PTR_BITWIDTH'b00001100001,
        `W_POS_PTR_BITWIDTH'b00001100100,
        `W_POS_PTR_BITWIDTH'b00001100111,
        `W_POS_PTR_BITWIDTH'b00001101010,
        `W_POS_PTR_BITWIDTH'b00001101101,
        `W_POS_PTR_BITWIDTH'b00001110000,
        `W_POS_PTR_BITWIDTH'b00001110011,
        `W_POS_PTR_BITWIDTH'b00001110110,
        `W_POS_PTR_BITWIDTH'b00001111001,
        `W_POS_PTR_BITWIDTH'b00001111100,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010000010,
        `W_POS_PTR_BITWIDTH'b00010000010
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00010000110,
        `W_POS_PTR_BITWIDTH'b00010001001,
        `W_POS_PTR_BITWIDTH'b00010001010,
        `W_POS_PTR_BITWIDTH'b00010001100,
        `W_POS_PTR_BITWIDTH'b00010001111,
        `W_POS_PTR_BITWIDTH'b00010010001,
        `W_POS_PTR_BITWIDTH'b00010010100,
        `W_POS_PTR_BITWIDTH'b00010010111,
        `W_POS_PTR_BITWIDTH'b00010011010,
        `W_POS_PTR_BITWIDTH'b00010011100,
        `W_POS_PTR_BITWIDTH'b00010011111,
        `W_POS_PTR_BITWIDTH'b00010100010,
        `W_POS_PTR_BITWIDTH'b00010100101,
        `W_POS_PTR_BITWIDTH'b00010100110,
        `W_POS_PTR_BITWIDTH'b00010101000,
        `W_POS_PTR_BITWIDTH'b00010101001,
        `W_POS_PTR_BITWIDTH'b00010101100,
        `W_POS_PTR_BITWIDTH'b00010101111,
        `W_POS_PTR_BITWIDTH'b00010110010,
        `W_POS_PTR_BITWIDTH'b00010110101,
        `W_POS_PTR_BITWIDTH'b00010110110,
        `W_POS_PTR_BITWIDTH'b00010111001,
        `W_POS_PTR_BITWIDTH'b00010111100,
        `W_POS_PTR_BITWIDTH'b00010111100
    };

// w_all
