// w_pos_ptr
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000000010,
        `W_POS_PTR_BITWIDTH'b00000000100,
        `W_POS_PTR_BITWIDTH'b00000000110,
        `W_POS_PTR_BITWIDTH'b00000001000,
        `W_POS_PTR_BITWIDTH'b00000001010,
        `W_POS_PTR_BITWIDTH'b00000001101,
        `W_POS_PTR_BITWIDTH'b00000010000,
        `W_POS_PTR_BITWIDTH'b00000010011,
        `W_POS_PTR_BITWIDTH'b00000010110,
        `W_POS_PTR_BITWIDTH'b00000011001,
        `W_POS_PTR_BITWIDTH'b00000011100,
        `W_POS_PTR_BITWIDTH'b00000011110,
        `W_POS_PTR_BITWIDTH'b00000100000,
        `W_POS_PTR_BITWIDTH'b00000100011,
        `W_POS_PTR_BITWIDTH'b00000100110,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000101100,
        `W_POS_PTR_BITWIDTH'b00000101110,
        `W_POS_PTR_BITWIDTH'b00000110000,
        `W_POS_PTR_BITWIDTH'b00000110011,
        `W_POS_PTR_BITWIDTH'b00000110101,
        `W_POS_PTR_BITWIDTH'b00000111000,
        `W_POS_PTR_BITWIDTH'b00000111010,
        `W_POS_PTR_BITWIDTH'b00000111100,
        `W_POS_PTR_BITWIDTH'b00000111111,
        `W_POS_PTR_BITWIDTH'b00001000010,
        `W_POS_PTR_BITWIDTH'b00001000100,
        `W_POS_PTR_BITWIDTH'b00001000111,
        `W_POS_PTR_BITWIDTH'b00001001010,
        `W_POS_PTR_BITWIDTH'b00001001101,
        `W_POS_PTR_BITWIDTH'b00001001110,
        `W_POS_PTR_BITWIDTH'b00001010000,
        `W_POS_PTR_BITWIDTH'b00001010010,
        `W_POS_PTR_BITWIDTH'b00001010101,
        `W_POS_PTR_BITWIDTH'b00001011000,
        `W_POS_PTR_BITWIDTH'b00001011011,
        `W_POS_PTR_BITWIDTH'b00001011110,
        `W_POS_PTR_BITWIDTH'b00001100001,
        `W_POS_PTR_BITWIDTH'b00001100100,
        `W_POS_PTR_BITWIDTH'b00001100110,
        `W_POS_PTR_BITWIDTH'b00001101000,
        `W_POS_PTR_BITWIDTH'b00001101011,
        `W_POS_PTR_BITWIDTH'b00001101101,
        `W_POS_PTR_BITWIDTH'b00001110000,
        `W_POS_PTR_BITWIDTH'b00001110010,
        `W_POS_PTR_BITWIDTH'b00001110101,
        `W_POS_PTR_BITWIDTH'b00001110101
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00001111011,
        `W_POS_PTR_BITWIDTH'b00001111101,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010000010,
        `W_POS_PTR_BITWIDTH'b00010000101,
        `W_POS_PTR_BITWIDTH'b00010001000,
        `W_POS_PTR_BITWIDTH'b00010001011,
        `W_POS_PTR_BITWIDTH'b00010001110,
        `W_POS_PTR_BITWIDTH'b00010010001,
        `W_POS_PTR_BITWIDTH'b00010010100,
        `W_POS_PTR_BITWIDTH'b00010010111,
        `W_POS_PTR_BITWIDTH'b00010011001,
        `W_POS_PTR_BITWIDTH'b00010011100,
        `W_POS_PTR_BITWIDTH'b00010011111,
        `W_POS_PTR_BITWIDTH'b00010100010,
        `W_POS_PTR_BITWIDTH'b00010100101,
        `W_POS_PTR_BITWIDTH'b00010101000,
        `W_POS_PTR_BITWIDTH'b00010101011,
        `W_POS_PTR_BITWIDTH'b00010101110,
        `W_POS_PTR_BITWIDTH'b00010110000,
        `W_POS_PTR_BITWIDTH'b00010110010,
        `W_POS_PTR_BITWIDTH'b00010110101,
        `W_POS_PTR_BITWIDTH'b00010111000,
        `W_POS_PTR_BITWIDTH'b00010111010,
        `W_POS_PTR_BITWIDTH'b00010111101,
        `W_POS_PTR_BITWIDTH'b00011000000,
        `W_POS_PTR_BITWIDTH'b00011000011,
        `W_POS_PTR_BITWIDTH'b00011000110,
        `W_POS_PTR_BITWIDTH'b00011001001,
        `W_POS_PTR_BITWIDTH'b00011001100,
        `W_POS_PTR_BITWIDTH'b00011001110,
        `W_POS_PTR_BITWIDTH'b00011010000,
        `W_POS_PTR_BITWIDTH'b00011010010,
        `W_POS_PTR_BITWIDTH'b00011010011,
        `W_POS_PTR_BITWIDTH'b00011010110,
        `W_POS_PTR_BITWIDTH'b00011011001,
        `W_POS_PTR_BITWIDTH'b00011011100,
        `W_POS_PTR_BITWIDTH'b00011011111,
        `W_POS_PTR_BITWIDTH'b00011100010,
        `W_POS_PTR_BITWIDTH'b00011100101,
        `W_POS_PTR_BITWIDTH'b00011101000,
        `W_POS_PTR_BITWIDTH'b00011101011,
        `W_POS_PTR_BITWIDTH'b00011101110,
        `W_POS_PTR_BITWIDTH'b00011110000,
        `W_POS_PTR_BITWIDTH'b00011110010,
        `W_POS_PTR_BITWIDTH'b00011110101,
        `W_POS_PTR_BITWIDTH'b00011111000,
        `W_POS_PTR_BITWIDTH'b00011111000
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00011111101,
        `W_POS_PTR_BITWIDTH'b00100000000,
        `W_POS_PTR_BITWIDTH'b00100000010,
        `W_POS_PTR_BITWIDTH'b00100000101,
        `W_POS_PTR_BITWIDTH'b00100001000,
        `W_POS_PTR_BITWIDTH'b00100001001,
        `W_POS_PTR_BITWIDTH'b00100001100,
        `W_POS_PTR_BITWIDTH'b00100001111,
        `W_POS_PTR_BITWIDTH'b00100010010,
        `W_POS_PTR_BITWIDTH'b00100010101,
        `W_POS_PTR_BITWIDTH'b00100011000,
        `W_POS_PTR_BITWIDTH'b00100011011,
        `W_POS_PTR_BITWIDTH'b00100011110,
        `W_POS_PTR_BITWIDTH'b00100100000,
        `W_POS_PTR_BITWIDTH'b00100100011,
        `W_POS_PTR_BITWIDTH'b00100100110,
        `W_POS_PTR_BITWIDTH'b00100101000,
        `W_POS_PTR_BITWIDTH'b00100101011,
        `W_POS_PTR_BITWIDTH'b00100101110,
        `W_POS_PTR_BITWIDTH'b00100110000,
        `W_POS_PTR_BITWIDTH'b00100110011,
        `W_POS_PTR_BITWIDTH'b00100110110,
        `W_POS_PTR_BITWIDTH'b00100111000,
        `W_POS_PTR_BITWIDTH'b00100111010,
        `W_POS_PTR_BITWIDTH'b00100111101,
        `W_POS_PTR_BITWIDTH'b00101000000,
        `W_POS_PTR_BITWIDTH'b00101000011,
        `W_POS_PTR_BITWIDTH'b00101000110,
        `W_POS_PTR_BITWIDTH'b00101001001,
        `W_POS_PTR_BITWIDTH'b00101001100,
        `W_POS_PTR_BITWIDTH'b00101001111,
        `W_POS_PTR_BITWIDTH'b00101010000,
        `W_POS_PTR_BITWIDTH'b00101010001,
        `W_POS_PTR_BITWIDTH'b00101010010,
        `W_POS_PTR_BITWIDTH'b00101010100,
        `W_POS_PTR_BITWIDTH'b00101010111,
        `W_POS_PTR_BITWIDTH'b00101011010,
        `W_POS_PTR_BITWIDTH'b00101011101,
        `W_POS_PTR_BITWIDTH'b00101011111,
        `W_POS_PTR_BITWIDTH'b00101100010,
        `W_POS_PTR_BITWIDTH'b00101100100,
        `W_POS_PTR_BITWIDTH'b00101100111,
        `W_POS_PTR_BITWIDTH'b00101101010,
        `W_POS_PTR_BITWIDTH'b00101101100,
        `W_POS_PTR_BITWIDTH'b00101101110,
        `W_POS_PTR_BITWIDTH'b00101110001,
        `W_POS_PTR_BITWIDTH'b00101110100,
        `W_POS_PTR_BITWIDTH'b00101110100
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00000000000,
        `W_POS_PTR_BITWIDTH'b00000001010,
        `W_POS_PTR_BITWIDTH'b00000010001,
        `W_POS_PTR_BITWIDTH'b00000011001,
        `W_POS_PTR_BITWIDTH'b00000011111,
        `W_POS_PTR_BITWIDTH'b00000101001,
        `W_POS_PTR_BITWIDTH'b00000110001,
        `W_POS_PTR_BITWIDTH'b00000111001,
        `W_POS_PTR_BITWIDTH'b00001000101,
        `W_POS_PTR_BITWIDTH'b00001010001,
        `W_POS_PTR_BITWIDTH'b00001011110,
        `W_POS_PTR_BITWIDTH'b00001100110,
        `W_POS_PTR_BITWIDTH'b00001110100,
        `W_POS_PTR_BITWIDTH'b00001111111,
        `W_POS_PTR_BITWIDTH'b00010001001,
        `W_POS_PTR_BITWIDTH'b00010010100,
        `W_POS_PTR_BITWIDTH'b00010011011,
        `W_POS_PTR_BITWIDTH'b00010100101,
        `W_POS_PTR_BITWIDTH'b00010101110,
        `W_POS_PTR_BITWIDTH'b00010110101,
        `W_POS_PTR_BITWIDTH'b00010111110,
        `W_POS_PTR_BITWIDTH'b00011000100,
        `W_POS_PTR_BITWIDTH'b00011001101,
        `W_POS_PTR_BITWIDTH'b00011010110,
        `W_POS_PTR_BITWIDTH'b00011100000,
        `W_POS_PTR_BITWIDTH'b00011101011,
        `W_POS_PTR_BITWIDTH'b00011111000,
        `W_POS_PTR_BITWIDTH'b00100000110,
        `W_POS_PTR_BITWIDTH'b00100010000,
        `W_POS_PTR_BITWIDTH'b00100011001,
        `W_POS_PTR_BITWIDTH'b00100011110,
        `W_POS_PTR_BITWIDTH'b00100101001,
        `W_POS_PTR_BITWIDTH'b00100110111,
        `W_POS_PTR_BITWIDTH'b00101000000,
        `W_POS_PTR_BITWIDTH'b00101001010,
        `W_POS_PTR_BITWIDTH'b00101010100,
        `W_POS_PTR_BITWIDTH'b00101100001,
        `W_POS_PTR_BITWIDTH'b00101101101,
        `W_POS_PTR_BITWIDTH'b00101110111,
        `W_POS_PTR_BITWIDTH'b00110000011,
        `W_POS_PTR_BITWIDTH'b00110001101,
        `W_POS_PTR_BITWIDTH'b00110010110,
        `W_POS_PTR_BITWIDTH'b00110011110,
        `W_POS_PTR_BITWIDTH'b00110100101,
        `W_POS_PTR_BITWIDTH'b00110101111,
        `W_POS_PTR_BITWIDTH'b00110110110,
        `W_POS_PTR_BITWIDTH'b00111000011,
        `W_POS_PTR_BITWIDTH'b00111000011
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
    '{
        `W_POS_PTR_BITWIDTH'b00111011010,
        `W_POS_PTR_BITWIDTH'b00111100100,
        `W_POS_PTR_BITWIDTH'b00111101110,
        `W_POS_PTR_BITWIDTH'b00111110111,
        `W_POS_PTR_BITWIDTH'b01000000000,
        `W_POS_PTR_BITWIDTH'b01000001000,
        `W_POS_PTR_BITWIDTH'b01000001110,
        `W_POS_PTR_BITWIDTH'b01000011000,
        `W_POS_PTR_BITWIDTH'b01000011110,
        `W_POS_PTR_BITWIDTH'b01000101010,
        `W_POS_PTR_BITWIDTH'b01000110101,
        `W_POS_PTR_BITWIDTH'b01001000010,
        `W_POS_PTR_BITWIDTH'b01001001111,
        `W_POS_PTR_BITWIDTH'b01001011100,
        `W_POS_PTR_BITWIDTH'b01001100001,
        `W_POS_PTR_BITWIDTH'b01001101011,
        `W_POS_PTR_BITWIDTH'b01001110100,
        `W_POS_PTR_BITWIDTH'b01001111100,
        `W_POS_PTR_BITWIDTH'b01010000100,
        `W_POS_PTR_BITWIDTH'b01010001111,
        `W_POS_PTR_BITWIDTH'b01010010111,
        `W_POS_PTR_BITWIDTH'b01010011110,
        `W_POS_PTR_BITWIDTH'b01010101010,
        `W_POS_PTR_BITWIDTH'b01010110010,
        `W_POS_PTR_BITWIDTH'b01010111110,
        `W_POS_PTR_BITWIDTH'b01011001000,
        `W_POS_PTR_BITWIDTH'b01011010101,
        `W_POS_PTR_BITWIDTH'b01011100010,
        `W_POS_PTR_BITWIDTH'b01011100111,
        `W_POS_PTR_BITWIDTH'b01011101111,
        `W_POS_PTR_BITWIDTH'b01011110100,
        `W_POS_PTR_BITWIDTH'b01100000000,
        `W_POS_PTR_BITWIDTH'b01100001000,
        `W_POS_PTR_BITWIDTH'b01100010001,
        `W_POS_PTR_BITWIDTH'b01100011011,
        `W_POS_PTR_BITWIDTH'b01100100101,
        `W_POS_PTR_BITWIDTH'b01100110100,
        `W_POS_PTR_BITWIDTH'b01100111111,
        `W_POS_PTR_BITWIDTH'b01101001000,
        `W_POS_PTR_BITWIDTH'b01101010011,
        `W_POS_PTR_BITWIDTH'b01101011111,
        `W_POS_PTR_BITWIDTH'b01101100111,
        `W_POS_PTR_BITWIDTH'b01101101101,
        `W_POS_PTR_BITWIDTH'b01101110111,
        `W_POS_PTR_BITWIDTH'b01101111110,
        `W_POS_PTR_BITWIDTH'b01110000101,
        `W_POS_PTR_BITWIDTH'b01110010001,
        `W_POS_PTR_BITWIDTH'b01110010001
    };
    localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
    '{
        `W_POS_PTR_BITWIDTH'b01110100110,
        `W_POS_PTR_BITWIDTH'b01110101100,
        `W_POS_PTR_BITWIDTH'b01110110011,
        `W_POS_PTR_BITWIDTH'b01110111011,
        `W_POS_PTR_BITWIDTH'b01111000011,
        `W_POS_PTR_BITWIDTH'b01111001011,
        `W_POS_PTR_BITWIDTH'b01111010010,
        `W_POS_PTR_BITWIDTH'b01111011110,
        `W_POS_PTR_BITWIDTH'b01111100111,
        `W_POS_PTR_BITWIDTH'b01111110001,
        `W_POS_PTR_BITWIDTH'b01111111101,
        `W_POS_PTR_BITWIDTH'b10000001001,
        `W_POS_PTR_BITWIDTH'b10000010101,
        `W_POS_PTR_BITWIDTH'b10000011111,
        `W_POS_PTR_BITWIDTH'b10000100111,
        `W_POS_PTR_BITWIDTH'b10000110100,
        `W_POS_PTR_BITWIDTH'b10000111100,
        `W_POS_PTR_BITWIDTH'b10001000110,
        `W_POS_PTR_BITWIDTH'b10001001110,
        `W_POS_PTR_BITWIDTH'b10001010100,
        `W_POS_PTR_BITWIDTH'b10001100001,
        `W_POS_PTR_BITWIDTH'b10001101100,
        `W_POS_PTR_BITWIDTH'b10001110111,
        `W_POS_PTR_BITWIDTH'b10010000000,
        `W_POS_PTR_BITWIDTH'b10010000110,
        `W_POS_PTR_BITWIDTH'b10010010001,
        `W_POS_PTR_BITWIDTH'b10010011011,
        `W_POS_PTR_BITWIDTH'b10010101001,
        `W_POS_PTR_BITWIDTH'b10010110010,
        `W_POS_PTR_BITWIDTH'b10010111000,
        `W_POS_PTR_BITWIDTH'b10011000000,
        `W_POS_PTR_BITWIDTH'b10011001011,
        `W_POS_PTR_BITWIDTH'b10011010100,
        `W_POS_PTR_BITWIDTH'b10011011100,
        `W_POS_PTR_BITWIDTH'b10011101100,
        `W_POS_PTR_BITWIDTH'b10011110111,
        `W_POS_PTR_BITWIDTH'b10100000011,
        `W_POS_PTR_BITWIDTH'b10100001100,
        `W_POS_PTR_BITWIDTH'b10100010101,
        `W_POS_PTR_BITWIDTH'b10100011110,
        `W_POS_PTR_BITWIDTH'b10100100011,
        `W_POS_PTR_BITWIDTH'b10100101100,
        `W_POS_PTR_BITWIDTH'b10100110100,
        `W_POS_PTR_BITWIDTH'b10100111011,
        `W_POS_PTR_BITWIDTH'b10100111111,
        `W_POS_PTR_BITWIDTH'b10101000001,
        `W_POS_PTR_BITWIDTH'b10101001101,
        `W_POS_PTR_BITWIDTH'b10101001101
    };

// w_pos_ptr
