`define W_DATA_BITWIDTH    16
`define W_C_BITWIDTH       5   // log2(# Channel)
`define W_R_BITWIDTH       2 
`define W_K_BITWIDTH       5 
`define W_POS_PTR_BITWIDTH 11 
// `define W_S_BITWIDTH       2  
// `define W_ITERS_BITWIDTH   6 


`define W_C_LENGTH_L1_S0  123
`define W_R_LENGTH_L1_S0  48
`define W_C_LENGTH_L1_S1  130
`define W_R_LENGTH_L1_S1  48
`define W_C_LENGTH_L1_S2  124
`define W_R_LENGTH_L1_S2  48

`define W_C_LENGTH_L2_S0  474
`define W_R_LENGTH_L2_S0  48
`define W_C_LENGTH_L2_S1  460
`define W_R_LENGTH_L2_S1  48
`define W_C_LENGTH_L2_S2  446
`define W_R_LENGTH_L2_S2  48

`define W_C_LENGTH_L3_S0  1136
`define W_R_LENGTH_L3_S0  96
`define W_C_LENGTH_L3_S1  1117
`define W_R_LENGTH_L3_S1  96
`define W_C_LENGTH_L3_S2  1131
`define W_R_LENGTH_L3_S2  96



module WMEM(
    input i_rst_n,
    input i_clk,
    // input i_start,
    // output logic o_finished,

    // w_data
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l3_s0 [0:`W_C_LENGTH_L3_S0-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l3_s1 [0:`W_C_LENGTH_L3_S1-1],
    output logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l3_s2 [0:`W_C_LENGTH_L3_S2-1],

    // w_c_idx
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l1_s0 [0:`W_C_LENGTH_L1_S0-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l1_s1 [0:`W_C_LENGTH_L1_S1-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l1_s2 [0:`W_C_LENGTH_L1_S2-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l2_s0 [0:`W_C_LENGTH_L2_S0-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l2_s1 [0:`W_C_LENGTH_L2_S1-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l2_s2 [0:`W_C_LENGTH_L2_S2-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l3_s0 [0:`W_C_LENGTH_L3_S0-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l3_s1 [0:`W_C_LENGTH_L3_S1-1],
    output logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l3_s2 [0:`W_C_LENGTH_L3_S2-1],

    // w_r_idx
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l3_s0 [0:`W_R_LENGTH_L3_S0-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l3_s1 [0:`W_R_LENGTH_L3_S1-1],
    output logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l3_s2 [0:`W_R_LENGTH_L3_S2-1],

    //  w_k_idx
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l3_s0 [0:`W_R_LENGTH_L3_S0-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l3_s1 [0:`W_R_LENGTH_L3_S1-1],
    output logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l3_s2 [0:`W_R_LENGTH_L3_S2-1],

    // w_pos_ptr
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l3_s0 [0:`W_R_LENGTH_L3_S0-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l3_s1 [0:`W_R_LENGTH_L3_S1-1],
    output logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l3_s2 [0:`W_R_LENGTH_L3_S2-1]
);

// ===== Parameters definition ===== 

// w_data
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
    '{
        `W_DATA_BITWIDTH'b11111_11101100110,
        `W_DATA_BITWIDTH'b11111_10111110001,
        `W_DATA_BITWIDTH'b00000_00010111001,
        `W_DATA_BITWIDTH'b11111_11001001000,
        `W_DATA_BITWIDTH'b11111_11100101100,
        `W_DATA_BITWIDTH'b11111_11101011010,
        `W_DATA_BITWIDTH'b00000_01011101001,
        `W_DATA_BITWIDTH'b00000_01110000101,
        `W_DATA_BITWIDTH'b11111_00101001100,
        `W_DATA_BITWIDTH'b11111_01000011010,
        `W_DATA_BITWIDTH'b00000_01000111111,
        `W_DATA_BITWIDTH'b11110_11110101000,
        `W_DATA_BITWIDTH'b11111_11011101100,
        `W_DATA_BITWIDTH'b00001_10100100001,
        `W_DATA_BITWIDTH'b00000_11110000000,
        `W_DATA_BITWIDTH'b11110_11101111100,
        `W_DATA_BITWIDTH'b00001_01111111011,
        `W_DATA_BITWIDTH'b11111_10110101010,
        `W_DATA_BITWIDTH'b00000_10000001010,
        `W_DATA_BITWIDTH'b00000_00010111010,
        `W_DATA_BITWIDTH'b11110_01101110010,
        `W_DATA_BITWIDTH'b00001_01101101000,
        `W_DATA_BITWIDTH'b00000_01101100100,
        `W_DATA_BITWIDTH'b00001_00001011110,
        `W_DATA_BITWIDTH'b11111_01101101010,
        `W_DATA_BITWIDTH'b00000_10110010101,
        `W_DATA_BITWIDTH'b00001_00011000111,
        `W_DATA_BITWIDTH'b11111_11001000000,
        `W_DATA_BITWIDTH'b11111_01000010001,
        `W_DATA_BITWIDTH'b00000_00111110100,
        `W_DATA_BITWIDTH'b00000_01111001101,
        `W_DATA_BITWIDTH'b00001_00001011110,
        `W_DATA_BITWIDTH'b00000_10110100100,
        `W_DATA_BITWIDTH'b00000_01001101110,
        `W_DATA_BITWIDTH'b11111_10000000001,
        `W_DATA_BITWIDTH'b11111_00111111011,
        `W_DATA_BITWIDTH'b11111_01010101100,
        `W_DATA_BITWIDTH'b11110_11110100100,
        `W_DATA_BITWIDTH'b00000_11011011001,
        `W_DATA_BITWIDTH'b11111_01111111110,
        `W_DATA_BITWIDTH'b00000_10000110000,
        `W_DATA_BITWIDTH'b11111_10110111010,
        `W_DATA_BITWIDTH'b11111_00011101101,
        `W_DATA_BITWIDTH'b11111_10010001101,
        `W_DATA_BITWIDTH'b00000_01110100011,
        `W_DATA_BITWIDTH'b00000_11111010101,
        `W_DATA_BITWIDTH'b11111_01110111101,
        `W_DATA_BITWIDTH'b00000_10101111100,
        `W_DATA_BITWIDTH'b00000_01011110110,
        `W_DATA_BITWIDTH'b00000_10010100011,
        `W_DATA_BITWIDTH'b00000_00100100010,
        `W_DATA_BITWIDTH'b00000_10110111000,
        `W_DATA_BITWIDTH'b00000_00100101001,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b00000_00111000001,
        `W_DATA_BITWIDTH'b11111_11100011101,
        `W_DATA_BITWIDTH'b11111_11001101111,
        `W_DATA_BITWIDTH'b11111_11000010110,
        `W_DATA_BITWIDTH'b00000_00111101010,
        `W_DATA_BITWIDTH'b00000_00111001111,
        `W_DATA_BITWIDTH'b11111_10101100100,
        `W_DATA_BITWIDTH'b00000_10001001100,
        `W_DATA_BITWIDTH'b00000_10010000011,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b00000_00100101011,
        `W_DATA_BITWIDTH'b00000_01001100011,
        `W_DATA_BITWIDTH'b11111_01111010111,
        `W_DATA_BITWIDTH'b11111_01010110111,
        `W_DATA_BITWIDTH'b00000_01111100111,
        `W_DATA_BITWIDTH'b00000_01101000010,
        `W_DATA_BITWIDTH'b11111_01110111001,
        `W_DATA_BITWIDTH'b00000_10010101110,
        `W_DATA_BITWIDTH'b00000_01111100110,
        `W_DATA_BITWIDTH'b00000_10010010110,
        `W_DATA_BITWIDTH'b11111_10100101101,
        `W_DATA_BITWIDTH'b11111_11011010101,
        `W_DATA_BITWIDTH'b11111_10100001000,
        `W_DATA_BITWIDTH'b11111_11011001011,
        `W_DATA_BITWIDTH'b11111_11100001010,
        `W_DATA_BITWIDTH'b11111_11010100111,
        `W_DATA_BITWIDTH'b11111_11001011111,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b11111_10101010000,
        `W_DATA_BITWIDTH'b11111_11001001110,
        `W_DATA_BITWIDTH'b11111_01010011110,
        `W_DATA_BITWIDTH'b11111_00100101111,
        `W_DATA_BITWIDTH'b11111_10010101000,
        `W_DATA_BITWIDTH'b11110_10110111011,
        `W_DATA_BITWIDTH'b00000_01011110000,
        `W_DATA_BITWIDTH'b11111_10010011011,
        `W_DATA_BITWIDTH'b00000_00111101001,
        `W_DATA_BITWIDTH'b00000_01101010010,
        `W_DATA_BITWIDTH'b00000_00010011101,
        `W_DATA_BITWIDTH'b11111_11000010111,
        `W_DATA_BITWIDTH'b00000_11110111111,
        `W_DATA_BITWIDTH'b00001_00010111000,
        `W_DATA_BITWIDTH'b00000_01000011010,
        `W_DATA_BITWIDTH'b11111_00110001010,
        `W_DATA_BITWIDTH'b11111_10011110100,
        `W_DATA_BITWIDTH'b11111_01011111011,
        `W_DATA_BITWIDTH'b00000_01011001011,
        `W_DATA_BITWIDTH'b00000_01000110010,
        `W_DATA_BITWIDTH'b11111_10010001011,
        `W_DATA_BITWIDTH'b11111_11101010100,
        `W_DATA_BITWIDTH'b11111_11101111110,
        `W_DATA_BITWIDTH'b00000_01001111101,
        `W_DATA_BITWIDTH'b00000_01000001111,
        `W_DATA_BITWIDTH'b11111_10111000001,
        `W_DATA_BITWIDTH'b11111_01000000010,
        `W_DATA_BITWIDTH'b00000_10000001111,
        `W_DATA_BITWIDTH'b11111_10101010001,
        `W_DATA_BITWIDTH'b00000_00101110110,
        `W_DATA_BITWIDTH'b00000_01100010100,
        `W_DATA_BITWIDTH'b00000_00011101010,
        `W_DATA_BITWIDTH'b00000_00110000101,
        `W_DATA_BITWIDTH'b11111_11100111100,
        `W_DATA_BITWIDTH'b00000_01000011100,
        `W_DATA_BITWIDTH'b00000_01000110011,
        `W_DATA_BITWIDTH'b00000_00110011001,
        `W_DATA_BITWIDTH'b00000_00101111100,
        `W_DATA_BITWIDTH'b00000_01001100000,
        `W_DATA_BITWIDTH'b11111_10110110110,
        `W_DATA_BITWIDTH'b11111_10110110110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
    '{
        `W_DATA_BITWIDTH'b00000_00101011111,
        `W_DATA_BITWIDTH'b00000_00010101011,
        `W_DATA_BITWIDTH'b00000_00111100111,
        `W_DATA_BITWIDTH'b00000_00100101110,
        `W_DATA_BITWIDTH'b00000_01000110010,
        `W_DATA_BITWIDTH'b11111_11010111000,
        `W_DATA_BITWIDTH'b11111_10111110110,
        `W_DATA_BITWIDTH'b11111_00111000001,
        `W_DATA_BITWIDTH'b11111_10111010101,
        `W_DATA_BITWIDTH'b11111_10000111010,
        `W_DATA_BITWIDTH'b00000_00100010000,
        `W_DATA_BITWIDTH'b00000_00011011000,
        `W_DATA_BITWIDTH'b11111_11010010100,
        `W_DATA_BITWIDTH'b00000_00101001111,
        `W_DATA_BITWIDTH'b11111_01100011101,
        `W_DATA_BITWIDTH'b00000_10110011010,
        `W_DATA_BITWIDTH'b11111_10100111010,
        `W_DATA_BITWIDTH'b11111_00010111110,
        `W_DATA_BITWIDTH'b11110_11101011101,
        `W_DATA_BITWIDTH'b11110_11000001011,
        `W_DATA_BITWIDTH'b11111_10101001011,
        `W_DATA_BITWIDTH'b00000_10111101111,
        `W_DATA_BITWIDTH'b11111_11000000100,
        `W_DATA_BITWIDTH'b00001_01110010000,
        `W_DATA_BITWIDTH'b11110_11100111010,
        `W_DATA_BITWIDTH'b00000_01101111000,
        `W_DATA_BITWIDTH'b11111_01010101101,
        `W_DATA_BITWIDTH'b00001_00000101000,
        `W_DATA_BITWIDTH'b00001_01110110101,
        `W_DATA_BITWIDTH'b11111_01100111000,
        `W_DATA_BITWIDTH'b11111_01100011100,
        `W_DATA_BITWIDTH'b11110_11100100010,
        `W_DATA_BITWIDTH'b00001_00000110000,
        `W_DATA_BITWIDTH'b00000_11110000000,
        `W_DATA_BITWIDTH'b00000_11000010101,
        `W_DATA_BITWIDTH'b00000_01010000011,
        `W_DATA_BITWIDTH'b00000_10000010000,
        `W_DATA_BITWIDTH'b00000_00011111110,
        `W_DATA_BITWIDTH'b11111_01100111110,
        `W_DATA_BITWIDTH'b11111_01110110110,
        `W_DATA_BITWIDTH'b00000_01000100110,
        `W_DATA_BITWIDTH'b00000_10011101111,
        `W_DATA_BITWIDTH'b00000_01010110001,
        `W_DATA_BITWIDTH'b00000_00010001101,
        `W_DATA_BITWIDTH'b11111_00011110100,
        `W_DATA_BITWIDTH'b11111_00110101001,
        `W_DATA_BITWIDTH'b00000_11101011110,
        `W_DATA_BITWIDTH'b11111_11011101000,
        `W_DATA_BITWIDTH'b00000_01110110001,
        `W_DATA_BITWIDTH'b00000_01101001111,
        `W_DATA_BITWIDTH'b00000_01110100111,
        `W_DATA_BITWIDTH'b11111_11011111010,
        `W_DATA_BITWIDTH'b11111_01000011110,
        `W_DATA_BITWIDTH'b11111_00110000110,
        `W_DATA_BITWIDTH'b00000_00111110100,
        `W_DATA_BITWIDTH'b11111_01011101001,
        `W_DATA_BITWIDTH'b11111_11011010000,
        `W_DATA_BITWIDTH'b00000_11100111011,
        `W_DATA_BITWIDTH'b11111_11001010001,
        `W_DATA_BITWIDTH'b00000_00011000101,
        `W_DATA_BITWIDTH'b00000_00100001001,
        `W_DATA_BITWIDTH'b11111_11101101011,
        `W_DATA_BITWIDTH'b11111_11010010000,
        `W_DATA_BITWIDTH'b00000_00010000011,
        `W_DATA_BITWIDTH'b00000_00110101011,
        `W_DATA_BITWIDTH'b00000_00011001110,
        `W_DATA_BITWIDTH'b00000_01011100010,
        `W_DATA_BITWIDTH'b11111_11001100000,
        `W_DATA_BITWIDTH'b00000_10000010010,
        `W_DATA_BITWIDTH'b00000_00100000100,
        `W_DATA_BITWIDTH'b11111_11011101001,
        `W_DATA_BITWIDTH'b11111_01101101001,
        `W_DATA_BITWIDTH'b11111_11101110000,
        `W_DATA_BITWIDTH'b11111_11100100110,
        `W_DATA_BITWIDTH'b11111_10011011001,
        `W_DATA_BITWIDTH'b11111_10011110101,
        `W_DATA_BITWIDTH'b00000_00110111011,
        `W_DATA_BITWIDTH'b00000_01000110011,
        `W_DATA_BITWIDTH'b11111_11010110001,
        `W_DATA_BITWIDTH'b00000_10010110111,
        `W_DATA_BITWIDTH'b00000_01000010010,
        `W_DATA_BITWIDTH'b00000_01111100010,
        `W_DATA_BITWIDTH'b11111_01110000101,
        `W_DATA_BITWIDTH'b11111_11100101011,
        `W_DATA_BITWIDTH'b00000_00010111010,
        `W_DATA_BITWIDTH'b11111_11100011011,
        `W_DATA_BITWIDTH'b00000_00100011110,
        `W_DATA_BITWIDTH'b11111_11101111001,
        `W_DATA_BITWIDTH'b11111_01111111100,
        `W_DATA_BITWIDTH'b00001_00011111111,
        `W_DATA_BITWIDTH'b00000_01001011111,
        `W_DATA_BITWIDTH'b11110_11100110011,
        `W_DATA_BITWIDTH'b00000_00101111010,
        `W_DATA_BITWIDTH'b00001_00001010011,
        `W_DATA_BITWIDTH'b00001_00100011011,
        `W_DATA_BITWIDTH'b11111_00011111100,
        `W_DATA_BITWIDTH'b00000_00011100010,
        `W_DATA_BITWIDTH'b00000_00110001010,
        `W_DATA_BITWIDTH'b00000_00101101101,
        `W_DATA_BITWIDTH'b00000_00100110111,
        `W_DATA_BITWIDTH'b11111_10000110011,
        `W_DATA_BITWIDTH'b11111_10011001100,
        `W_DATA_BITWIDTH'b00000_10011110100,
        `W_DATA_BITWIDTH'b11111_00001111001,
        `W_DATA_BITWIDTH'b11111_01011000000,
        `W_DATA_BITWIDTH'b00000_11000110100,
        `W_DATA_BITWIDTH'b11111_11000010010,
        `W_DATA_BITWIDTH'b11111_10101110110,
        `W_DATA_BITWIDTH'b11111_10000001110,
        `W_DATA_BITWIDTH'b11111_10101100100,
        `W_DATA_BITWIDTH'b00000_01110111111,
        `W_DATA_BITWIDTH'b11111_11101110011,
        `W_DATA_BITWIDTH'b00000_00111101110,
        `W_DATA_BITWIDTH'b00000_01100100011,
        `W_DATA_BITWIDTH'b11111_10110110100,
        `W_DATA_BITWIDTH'b11111_11100110101,
        `W_DATA_BITWIDTH'b00000_00111111110,
        `W_DATA_BITWIDTH'b00000_01101111010,
        `W_DATA_BITWIDTH'b11111_11000111010,
        `W_DATA_BITWIDTH'b11111_11101010101,
        `W_DATA_BITWIDTH'b11111_10010000001,
        `W_DATA_BITWIDTH'b11111_10000111011,
        `W_DATA_BITWIDTH'b11111_10110111010,
        `W_DATA_BITWIDTH'b11111_11001000010,
        `W_DATA_BITWIDTH'b11111_11001101010,
        `W_DATA_BITWIDTH'b11111_10111110111,
        `W_DATA_BITWIDTH'b00000_00111000111,
        `W_DATA_BITWIDTH'b00000_01011100000,
        `W_DATA_BITWIDTH'b00000_00101101011,
        `W_DATA_BITWIDTH'b00000_00101101011
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
    '{
        `W_DATA_BITWIDTH'b00000_00011001100,
        `W_DATA_BITWIDTH'b11111_11001101101,
        `W_DATA_BITWIDTH'b00000_00011011100,
        `W_DATA_BITWIDTH'b00000_00101101111,
        `W_DATA_BITWIDTH'b00000_00011000011,
        `W_DATA_BITWIDTH'b00000_00110001110,
        `W_DATA_BITWIDTH'b00000_00111000011,
        `W_DATA_BITWIDTH'b00000_00100111000,
        `W_DATA_BITWIDTH'b00000_01010100011,
        `W_DATA_BITWIDTH'b00000_11001010111,
        `W_DATA_BITWIDTH'b00000_10111100000,
        `W_DATA_BITWIDTH'b11111_10101010110,
        `W_DATA_BITWIDTH'b00000_01110110110,
        `W_DATA_BITWIDTH'b00000_10000001100,
        `W_DATA_BITWIDTH'b00000_11101011110,
        `W_DATA_BITWIDTH'b00001_00011000010,
        `W_DATA_BITWIDTH'b00000_00100011101,
        `W_DATA_BITWIDTH'b00000_10110101000,
        `W_DATA_BITWIDTH'b11111_10111000001,
        `W_DATA_BITWIDTH'b11111_01101110010,
        `W_DATA_BITWIDTH'b11111_00001100100,
        `W_DATA_BITWIDTH'b11110_11100010000,
        `W_DATA_BITWIDTH'b00000_01010010010,
        `W_DATA_BITWIDTH'b00001_00010011111,
        `W_DATA_BITWIDTH'b11111_11001101100,
        `W_DATA_BITWIDTH'b11111_00000100001,
        `W_DATA_BITWIDTH'b11111_10001100011,
        `W_DATA_BITWIDTH'b11111_10101110110,
        `W_DATA_BITWIDTH'b00000_00010100111,
        `W_DATA_BITWIDTH'b11110_11101000001,
        `W_DATA_BITWIDTH'b11110_11110011101,
        `W_DATA_BITWIDTH'b00000_00100001110,
        `W_DATA_BITWIDTH'b00000_01110110100,
        `W_DATA_BITWIDTH'b11111_01101011100,
        `W_DATA_BITWIDTH'b00000_00110010011,
        `W_DATA_BITWIDTH'b11111_01000101111,
        `W_DATA_BITWIDTH'b11111_11001100001,
        `W_DATA_BITWIDTH'b11111_10000101001,
        `W_DATA_BITWIDTH'b11111_01101110000,
        `W_DATA_BITWIDTH'b00000_01101010011,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b00000_10011110101,
        `W_DATA_BITWIDTH'b11111_00010100000,
        `W_DATA_BITWIDTH'b11110_11000000110,
        `W_DATA_BITWIDTH'b11111_01001101111,
        `W_DATA_BITWIDTH'b11111_10101000000,
        `W_DATA_BITWIDTH'b00000_01011000000,
        `W_DATA_BITWIDTH'b00000_11010001000,
        `W_DATA_BITWIDTH'b00000_01000110001,
        `W_DATA_BITWIDTH'b00000_10111001000,
        `W_DATA_BITWIDTH'b11111_01010011000,
        `W_DATA_BITWIDTH'b11111_00001101011,
        `W_DATA_BITWIDTH'b11111_11011001100,
        `W_DATA_BITWIDTH'b11111_00010111100,
        `W_DATA_BITWIDTH'b00000_01110101000,
        `W_DATA_BITWIDTH'b00000_00100011011,
        `W_DATA_BITWIDTH'b00000_11111001100,
        `W_DATA_BITWIDTH'b00000_00010101000,
        `W_DATA_BITWIDTH'b00000_00100111010,
        `W_DATA_BITWIDTH'b00000_00101100011,
        `W_DATA_BITWIDTH'b11111_11011001101,
        `W_DATA_BITWIDTH'b00000_01001000110,
        `W_DATA_BITWIDTH'b00000_01001000011,
        `W_DATA_BITWIDTH'b11111_11011101110,
        `W_DATA_BITWIDTH'b00000_01110000101,
        `W_DATA_BITWIDTH'b00000_01110011101,
        `W_DATA_BITWIDTH'b11111_11000001111,
        `W_DATA_BITWIDTH'b00000_01011110001,
        `W_DATA_BITWIDTH'b00000_00010111010,
        `W_DATA_BITWIDTH'b00000_00100100001,
        `W_DATA_BITWIDTH'b00000_01011111111,
        `W_DATA_BITWIDTH'b11111_10101010110,
        `W_DATA_BITWIDTH'b11111_11011100001,
        `W_DATA_BITWIDTH'b11111_01101010001,
        `W_DATA_BITWIDTH'b11111_10001110111,
        `W_DATA_BITWIDTH'b00000_01010111101,
        `W_DATA_BITWIDTH'b11111_10001101001,
        `W_DATA_BITWIDTH'b00000_01010100110,
        `W_DATA_BITWIDTH'b00000_01101010001,
        `W_DATA_BITWIDTH'b11111_10001001111,
        `W_DATA_BITWIDTH'b11111_11010101010,
        `W_DATA_BITWIDTH'b11111_11011100110,
        `W_DATA_BITWIDTH'b00000_00100001110,
        `W_DATA_BITWIDTH'b00000_00101000111,
        `W_DATA_BITWIDTH'b11111_11011110011,
        `W_DATA_BITWIDTH'b00000_10111010101,
        `W_DATA_BITWIDTH'b00000_11011111100,
        `W_DATA_BITWIDTH'b00000_11010010110,
        `W_DATA_BITWIDTH'b00000_01000100010,
        `W_DATA_BITWIDTH'b11111_01010000010,
        `W_DATA_BITWIDTH'b11111_11000101001,
        `W_DATA_BITWIDTH'b11111_10110010100,
        `W_DATA_BITWIDTH'b00000_00111011110,
        `W_DATA_BITWIDTH'b11111_01011011110,
        `W_DATA_BITWIDTH'b00000_11111111101,
        `W_DATA_BITWIDTH'b11110_11101110110,
        `W_DATA_BITWIDTH'b11111_10111011101,
        `W_DATA_BITWIDTH'b11111_11000101110,
        `W_DATA_BITWIDTH'b00000_10011001111,
        `W_DATA_BITWIDTH'b00000_01010011000,
        `W_DATA_BITWIDTH'b11111_01011100110,
        `W_DATA_BITWIDTH'b11111_11000011100,
        `W_DATA_BITWIDTH'b11111_11000010110,
        `W_DATA_BITWIDTH'b11111_10101011010,
        `W_DATA_BITWIDTH'b11111_10101001001,
        `W_DATA_BITWIDTH'b11111_11001100010,
        `W_DATA_BITWIDTH'b00000_00110110101,
        `W_DATA_BITWIDTH'b00000_00110111010,
        `W_DATA_BITWIDTH'b00000_00010100111,
        `W_DATA_BITWIDTH'b00000_01011100010,
        `W_DATA_BITWIDTH'b00000_00010100110,
        `W_DATA_BITWIDTH'b00000_01010000000,
        `W_DATA_BITWIDTH'b11111_11001011011,
        `W_DATA_BITWIDTH'b11111_11011011111,
        `W_DATA_BITWIDTH'b11111_10001101000,
        `W_DATA_BITWIDTH'b11111_10111010101,
        `W_DATA_BITWIDTH'b11111_11010100010,
        `W_DATA_BITWIDTH'b11111_11001011001,
        `W_DATA_BITWIDTH'b11111_11001111110,
        `W_DATA_BITWIDTH'b00000_01010101001,
        `W_DATA_BITWIDTH'b11111_11001011110,
        `W_DATA_BITWIDTH'b00000_00100010001,
        `W_DATA_BITWIDTH'b11111_11000010110,
        `W_DATA_BITWIDTH'b11111_11000010110
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
    '{
        `W_DATA_BITWIDTH'b00000_00010101111,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b00000_00011111100,
        `W_DATA_BITWIDTH'b11111_11011001111,
        `W_DATA_BITWIDTH'b11111_11101110101,
        `W_DATA_BITWIDTH'b11111_11101101010,
        `W_DATA_BITWIDTH'b11111_11100001010,
        `W_DATA_BITWIDTH'b11111_11001010010,
        `W_DATA_BITWIDTH'b11111_11100100111,
        `W_DATA_BITWIDTH'b11111_11101101011,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b00000_00010011110,
        `W_DATA_BITWIDTH'b00000_00010011110,
        `W_DATA_BITWIDTH'b11111_11101010111,
        `W_DATA_BITWIDTH'b00000_00010011101,
        `W_DATA_BITWIDTH'b11111_11011010101,
        `W_DATA_BITWIDTH'b00000_00011011001,
        `W_DATA_BITWIDTH'b00000_00100110100,
        `W_DATA_BITWIDTH'b11111_11100100000,
        `W_DATA_BITWIDTH'b00000_00010000011,
        `W_DATA_BITWIDTH'b00000_00010010010,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b00000_00110001101,
        `W_DATA_BITWIDTH'b11111_11010111110,
        `W_DATA_BITWIDTH'b00000_00010100111,
        `W_DATA_BITWIDTH'b11111_11101001111,
        `W_DATA_BITWIDTH'b00000_00101001001,
        `W_DATA_BITWIDTH'b00000_00010101111,
        `W_DATA_BITWIDTH'b00000_00010001000,
        `W_DATA_BITWIDTH'b11111_11101001110,
        `W_DATA_BITWIDTH'b11111_11100000100,
        `W_DATA_BITWIDTH'b00000_00010111100,
        `W_DATA_BITWIDTH'b00000_00011101000,
        `W_DATA_BITWIDTH'b11111_11101100111,
        `W_DATA_BITWIDTH'b00000_00010100001,
        `W_DATA_BITWIDTH'b11111_11011100111,
        `W_DATA_BITWIDTH'b11111_11101101001,
        `W_DATA_BITWIDTH'b00000_00010011111,
        `W_DATA_BITWIDTH'b11111_11100001000,
        `W_DATA_BITWIDTH'b00000_00011000010,
        `W_DATA_BITWIDTH'b00000_00010100100,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b00000_00011011100,
        `W_DATA_BITWIDTH'b00000_00010101101,
        `W_DATA_BITWIDTH'b11111_11100011011,
        `W_DATA_BITWIDTH'b11111_11011000111,
        `W_DATA_BITWIDTH'b00000_00011000000,
        `W_DATA_BITWIDTH'b00000_00011110111,
        `W_DATA_BITWIDTH'b00000_00010111101,
        `W_DATA_BITWIDTH'b11111_11011100100,
        `W_DATA_BITWIDTH'b11111_11001110100,
        `W_DATA_BITWIDTH'b11111_11001000101,
        `W_DATA_BITWIDTH'b00000_00100111001,
        `W_DATA_BITWIDTH'b11111_11100101011,
        `W_DATA_BITWIDTH'b00000_00110001111,
        `W_DATA_BITWIDTH'b11111_11101010111,
        `W_DATA_BITWIDTH'b00000_00101100010,
        `W_DATA_BITWIDTH'b11111_11100001101,
        `W_DATA_BITWIDTH'b00000_00010000010,
        `W_DATA_BITWIDTH'b11111_11011010110,
        `W_DATA_BITWIDTH'b00000_00011011101,
        `W_DATA_BITWIDTH'b11111_10111000000,
        `W_DATA_BITWIDTH'b11111_11001011011,
        `W_DATA_BITWIDTH'b11111_11000101101,
        `W_DATA_BITWIDTH'b00000_00100101110,
        `W_DATA_BITWIDTH'b00000_00011100011,
        `W_DATA_BITWIDTH'b11111_11100011101,
        `W_DATA_BITWIDTH'b11111_11101100011,
        `W_DATA_BITWIDTH'b11111_10111110011,
        `W_DATA_BITWIDTH'b11111_11010011010,
        `W_DATA_BITWIDTH'b00000_00010011000,
        `W_DATA_BITWIDTH'b11111_11101011101,
        `W_DATA_BITWIDTH'b00000_00100010011,
        `W_DATA_BITWIDTH'b11111_11011011000,
        `W_DATA_BITWIDTH'b11111_11101000011,
        `W_DATA_BITWIDTH'b11111_11101000110,
        `W_DATA_BITWIDTH'b00000_00100010110,
        `W_DATA_BITWIDTH'b00000_00011100001,
        `W_DATA_BITWIDTH'b11111_11011011010,
        `W_DATA_BITWIDTH'b11111_10111011001,
        `W_DATA_BITWIDTH'b11111_11010110110,
        `W_DATA_BITWIDTH'b11111_11011001010,
        `W_DATA_BITWIDTH'b00000_00100001011,
        `W_DATA_BITWIDTH'b00000_00010010100,
        `W_DATA_BITWIDTH'b11111_11011001110,
        `W_DATA_BITWIDTH'b11111_11001100010,
        `W_DATA_BITWIDTH'b00000_00010100101,
        `W_DATA_BITWIDTH'b11111_11010101110,
        `W_DATA_BITWIDTH'b11111_11101010101,
        `W_DATA_BITWIDTH'b11111_11010101000,
        `W_DATA_BITWIDTH'b11111_11100111001,
        `W_DATA_BITWIDTH'b11111_11010110010,
        `W_DATA_BITWIDTH'b00000_00010110101,
        `W_DATA_BITWIDTH'b11111_11100110100,
        `W_DATA_BITWIDTH'b11111_11100011100,
        `W_DATA_BITWIDTH'b11111_10110001010,
        `W_DATA_BITWIDTH'b00000_00010110111,
        `W_DATA_BITWIDTH'b00000_00111001000,
        `W_DATA_BITWIDTH'b00000_00100101101,
        `W_DATA_BITWIDTH'b11111_11010111001,
        `W_DATA_BITWIDTH'b00000_00011001101,
        `W_DATA_BITWIDTH'b11111_10001110111,
        `W_DATA_BITWIDTH'b11111_11000100001,
        `W_DATA_BITWIDTH'b00000_00100001111,
        `W_DATA_BITWIDTH'b11111_10100001001,
        `W_DATA_BITWIDTH'b11111_11010010111,
        `W_DATA_BITWIDTH'b11111_10111001110,
        `W_DATA_BITWIDTH'b00000_00011001100,
        `W_DATA_BITWIDTH'b11111_11001001100,
        `W_DATA_BITWIDTH'b11111_10110100001,
        `W_DATA_BITWIDTH'b11111_11011010010,
        `W_DATA_BITWIDTH'b00000_00101110000,
        `W_DATA_BITWIDTH'b11111_11010111010,
        `W_DATA_BITWIDTH'b11111_11011101010,
        `W_DATA_BITWIDTH'b11111_11010100011,
        `W_DATA_BITWIDTH'b11111_11101010111,
        `W_DATA_BITWIDTH'b11111_11100100101,
        `W_DATA_BITWIDTH'b11111_11100000010,
        `W_DATA_BITWIDTH'b11111_11011011011,
        `W_DATA_BITWIDTH'b00000_00100110100,
        `W_DATA_BITWIDTH'b11111_11100111011,
        `W_DATA_BITWIDTH'b00000_00011010111,
        `W_DATA_BITWIDTH'b11111_11100011011,
        `W_DATA_BITWIDTH'b11111_11101100000,
        `W_DATA_BITWIDTH'b00000_00010110010,
        `W_DATA_BITWIDTH'b11111_11100101101,
        `W_DATA_BITWIDTH'b00000_00100101110,
        `W_DATA_BITWIDTH'b00000_00010100000,
        `W_DATA_BITWIDTH'b11111_11010010101,
        `W_DATA_BITWIDTH'b11111_11101001100,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b11111_11010110101,
        `W_DATA_BITWIDTH'b11111_11101111100,
        `W_DATA_BITWIDTH'b00000_00010111111,
        `W_DATA_BITWIDTH'b11111_11010100100,
        `W_DATA_BITWIDTH'b00000_00011110111,
        `W_DATA_BITWIDTH'b11111_11100110111,
        `W_DATA_BITWIDTH'b11111_11011011100,
        `W_DATA_BITWIDTH'b11111_11100001011,
        `W_DATA_BITWIDTH'b11111_11100011101,
        `W_DATA_BITWIDTH'b11111_11100101110,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b11111_11101100111,
        `W_DATA_BITWIDTH'b11111_11011110000,
        `W_DATA_BITWIDTH'b11111_11100100000,
        `W_DATA_BITWIDTH'b00000_00100011111,
        `W_DATA_BITWIDTH'b00000_00100100101,
        `W_DATA_BITWIDTH'b11111_11100011000,
        `W_DATA_BITWIDTH'b11111_11010100010,
        `W_DATA_BITWIDTH'b11111_11010110000,
        `W_DATA_BITWIDTH'b00000_00010111011,
        `W_DATA_BITWIDTH'b00000_00010100001,
        `W_DATA_BITWIDTH'b11111_11001100110,
        `W_DATA_BITWIDTH'b00000_00010000100,
        `W_DATA_BITWIDTH'b00000_00011010000,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b00000_00010101011,
        `W_DATA_BITWIDTH'b00000_00011000010,
        `W_DATA_BITWIDTH'b00000_00100001101,
        `W_DATA_BITWIDTH'b00000_00011101101,
        `W_DATA_BITWIDTH'b00000_00010001101,
        `W_DATA_BITWIDTH'b11111_11101101011,
        `W_DATA_BITWIDTH'b11111_11011101101,
        `W_DATA_BITWIDTH'b11111_11101101000,
        `W_DATA_BITWIDTH'b11111_11101011110,
        `W_DATA_BITWIDTH'b00000_00100010111,
        `W_DATA_BITWIDTH'b11111_11100100011,
        `W_DATA_BITWIDTH'b00000_00101001001,
        `W_DATA_BITWIDTH'b00000_00011000000,
        `W_DATA_BITWIDTH'b00000_00101110110,
        `W_DATA_BITWIDTH'b00000_00010110110,
        `W_DATA_BITWIDTH'b11111_11101111010,
        `W_DATA_BITWIDTH'b00000_00100011101,
        `W_DATA_BITWIDTH'b00000_00011010011,
        `W_DATA_BITWIDTH'b00000_00010000110,
        `W_DATA_BITWIDTH'b11111_11100100010,
        `W_DATA_BITWIDTH'b11111_11011110011,
        `W_DATA_BITWIDTH'b00000_00010000001,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b00000_00011100001,
        `W_DATA_BITWIDTH'b00000_00011000011,
        `W_DATA_BITWIDTH'b11111_11101001001,
        `W_DATA_BITWIDTH'b11111_11101010001,
        `W_DATA_BITWIDTH'b11111_11101100101,
        `W_DATA_BITWIDTH'b11111_11100101111,
        `W_DATA_BITWIDTH'b11111_11100001011,
        `W_DATA_BITWIDTH'b00000_00011111100,
        `W_DATA_BITWIDTH'b11111_11100000010,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b00000_00011100011,
        `W_DATA_BITWIDTH'b11111_11100010000,
        `W_DATA_BITWIDTH'b11111_11010101110,
        `W_DATA_BITWIDTH'b11111_11011000011,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b11111_11011110101,
        `W_DATA_BITWIDTH'b11111_11011010011,
        `W_DATA_BITWIDTH'b11111_11101000000,
        `W_DATA_BITWIDTH'b11111_11001111100,
        `W_DATA_BITWIDTH'b11111_11001100110,
        `W_DATA_BITWIDTH'b00000_00011101000,
        `W_DATA_BITWIDTH'b11111_11101101111,
        `W_DATA_BITWIDTH'b00000_00010110001,
        `W_DATA_BITWIDTH'b00000_00011101010,
        `W_DATA_BITWIDTH'b11111_11101100110,
        `W_DATA_BITWIDTH'b00000_00010111001,
        `W_DATA_BITWIDTH'b11111_11101101011,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b00000_00100010010,
        `W_DATA_BITWIDTH'b00000_00100110100,
        `W_DATA_BITWIDTH'b00000_00010111111,
        `W_DATA_BITWIDTH'b11111_11010110110,
        `W_DATA_BITWIDTH'b11111_11100111110,
        `W_DATA_BITWIDTH'b00000_00100001010,
        `W_DATA_BITWIDTH'b11111_11101010000,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b11111_11101111001,
        `W_DATA_BITWIDTH'b00000_00101111001,
        `W_DATA_BITWIDTH'b00000_00010101110,
        `W_DATA_BITWIDTH'b11111_11011101110,
        `W_DATA_BITWIDTH'b00000_00101111101,
        `W_DATA_BITWIDTH'b11111_11100100111,
        `W_DATA_BITWIDTH'b00000_00010001011,
        `W_DATA_BITWIDTH'b00000_00011101010,
        `W_DATA_BITWIDTH'b11111_11010100011,
        `W_DATA_BITWIDTH'b00000_00100100011,
        `W_DATA_BITWIDTH'b00000_00010011110,
        `W_DATA_BITWIDTH'b11111_10110111010,
        `W_DATA_BITWIDTH'b11111_11101000110,
        `W_DATA_BITWIDTH'b11111_11011001000,
        `W_DATA_BITWIDTH'b00000_00011010001,
        `W_DATA_BITWIDTH'b11111_10001011000,
        `W_DATA_BITWIDTH'b11111_11100000100,
        `W_DATA_BITWIDTH'b00000_00111001101,
        `W_DATA_BITWIDTH'b11111_11100101000,
        `W_DATA_BITWIDTH'b00000_00101001011,
        `W_DATA_BITWIDTH'b00000_00110110111,
        `W_DATA_BITWIDTH'b11111_10101001010,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b00000_01000010101,
        `W_DATA_BITWIDTH'b11111_11001010010,
        `W_DATA_BITWIDTH'b00000_00110001000,
        `W_DATA_BITWIDTH'b00000_00011100110,
        `W_DATA_BITWIDTH'b11111_10111000110,
        `W_DATA_BITWIDTH'b11111_11001101001,
        `W_DATA_BITWIDTH'b11111_11001110011,
        `W_DATA_BITWIDTH'b11111_11101001010,
        `W_DATA_BITWIDTH'b11111_11011000000,
        `W_DATA_BITWIDTH'b00000_00101010010,
        `W_DATA_BITWIDTH'b00000_00100101000,
        `W_DATA_BITWIDTH'b11111_11010011010,
        `W_DATA_BITWIDTH'b11111_11001111100,
        `W_DATA_BITWIDTH'b11111_11100000011,
        `W_DATA_BITWIDTH'b00000_00011000111,
        `W_DATA_BITWIDTH'b00000_00110001101,
        `W_DATA_BITWIDTH'b11111_11101001011,
        `W_DATA_BITWIDTH'b11111_11010111110,
        `W_DATA_BITWIDTH'b11111_11001100101,
        `W_DATA_BITWIDTH'b00000_01000110111,
        `W_DATA_BITWIDTH'b11111_11000100010,
        `W_DATA_BITWIDTH'b11111_11100011001,
        `W_DATA_BITWIDTH'b00000_01001000111,
        `W_DATA_BITWIDTH'b00000_00100000101,
        `W_DATA_BITWIDTH'b00000_00011101110,
        `W_DATA_BITWIDTH'b11111_11100011101,
        `W_DATA_BITWIDTH'b11111_11101000101,
        `W_DATA_BITWIDTH'b11111_11101111100,
        `W_DATA_BITWIDTH'b11111_11100110100,
        `W_DATA_BITWIDTH'b11111_11100101010,
        `W_DATA_BITWIDTH'b00000_00010010100,
        `W_DATA_BITWIDTH'b11111_11100101010,
        `W_DATA_BITWIDTH'b11111_11101010010,
        `W_DATA_BITWIDTH'b11111_11011110001,
        `W_DATA_BITWIDTH'b11111_11001001011,
        `W_DATA_BITWIDTH'b00000_00011101110,
        `W_DATA_BITWIDTH'b11111_11101110000,
        `W_DATA_BITWIDTH'b11111_11101011100,
        `W_DATA_BITWIDTH'b11111_11100110100,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b00000_00100011111,
        `W_DATA_BITWIDTH'b11111_11100010100,
        `W_DATA_BITWIDTH'b11111_11101110111,
        `W_DATA_BITWIDTH'b00000_00010001100,
        `W_DATA_BITWIDTH'b11111_11011001110,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b00000_00100001101,
        `W_DATA_BITWIDTH'b11111_11100101011,
        `W_DATA_BITWIDTH'b11111_11101011100,
        `W_DATA_BITWIDTH'b00000_00101100010,
        `W_DATA_BITWIDTH'b00000_00011001001,
        `W_DATA_BITWIDTH'b11111_11011100101,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b00000_00011100010,
        `W_DATA_BITWIDTH'b00000_00100011100,
        `W_DATA_BITWIDTH'b11111_11011100111,
        `W_DATA_BITWIDTH'b00000_00110000011,
        `W_DATA_BITWIDTH'b11111_11100000000,
        `W_DATA_BITWIDTH'b11111_11011111010,
        `W_DATA_BITWIDTH'b00000_00100011101,
        `W_DATA_BITWIDTH'b11111_11011110010,
        `W_DATA_BITWIDTH'b11111_11100101110,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b11111_11000010001,
        `W_DATA_BITWIDTH'b11111_11101100110,
        `W_DATA_BITWIDTH'b11111_11010101010,
        `W_DATA_BITWIDTH'b11111_11011100100,
        `W_DATA_BITWIDTH'b11111_11011100000,
        `W_DATA_BITWIDTH'b11111_11100011000,
        `W_DATA_BITWIDTH'b11111_11100100100,
        `W_DATA_BITWIDTH'b11111_11101101110,
        `W_DATA_BITWIDTH'b11111_11101101100,
        `W_DATA_BITWIDTH'b00000_00010100011,
        `W_DATA_BITWIDTH'b11111_11001010001,
        `W_DATA_BITWIDTH'b11111_11101000010,
        `W_DATA_BITWIDTH'b11111_11011111100,
        `W_DATA_BITWIDTH'b11111_11010100100,
        `W_DATA_BITWIDTH'b11111_11010111111,
        `W_DATA_BITWIDTH'b00000_00010001010,
        `W_DATA_BITWIDTH'b11111_11100101000,
        `W_DATA_BITWIDTH'b11111_11000101010,
        `W_DATA_BITWIDTH'b00000_00100101101,
        `W_DATA_BITWIDTH'b00000_01001100010,
        `W_DATA_BITWIDTH'b11111_11100101111,
        `W_DATA_BITWIDTH'b11111_11100111000,
        `W_DATA_BITWIDTH'b11111_11101110111,
        `W_DATA_BITWIDTH'b00000_01010100001,
        `W_DATA_BITWIDTH'b00000_00011001010,
        `W_DATA_BITWIDTH'b00000_00010110001,
        `W_DATA_BITWIDTH'b00000_00011011100,
        `W_DATA_BITWIDTH'b11111_11011111010,
        `W_DATA_BITWIDTH'b11111_11100111111,
        `W_DATA_BITWIDTH'b00000_00110001110,
        `W_DATA_BITWIDTH'b11111_11100100001,
        `W_DATA_BITWIDTH'b11111_11100111000,
        `W_DATA_BITWIDTH'b11111_11010101101,
        `W_DATA_BITWIDTH'b00000_00100111010,
        `W_DATA_BITWIDTH'b11111_11100110110,
        `W_DATA_BITWIDTH'b00000_00100011010,
        `W_DATA_BITWIDTH'b11111_11100110011,
        `W_DATA_BITWIDTH'b00000_00110101000,
        `W_DATA_BITWIDTH'b00000_00011000000,
        `W_DATA_BITWIDTH'b00000_00111011000,
        `W_DATA_BITWIDTH'b00000_00010001100,
        `W_DATA_BITWIDTH'b00000_00111100110,
        `W_DATA_BITWIDTH'b11111_11011111101,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b00000_00110011101,
        `W_DATA_BITWIDTH'b11111_11101111011,
        `W_DATA_BITWIDTH'b11111_11000111001,
        `W_DATA_BITWIDTH'b11111_11001100110,
        `W_DATA_BITWIDTH'b11111_11001001001,
        `W_DATA_BITWIDTH'b00000_00111111000,
        `W_DATA_BITWIDTH'b11111_11001111011,
        `W_DATA_BITWIDTH'b00000_00011011100,
        `W_DATA_BITWIDTH'b11111_11011010010,
        `W_DATA_BITWIDTH'b11111_11000011001,
        `W_DATA_BITWIDTH'b00000_00010001010,
        `W_DATA_BITWIDTH'b11111_11101010101,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b11111_11010000011,
        `W_DATA_BITWIDTH'b00000_00011000110,
        `W_DATA_BITWIDTH'b11111_11001111010,
        `W_DATA_BITWIDTH'b11111_10111011001,
        `W_DATA_BITWIDTH'b11111_11101010001,
        `W_DATA_BITWIDTH'b11111_11001110011,
        `W_DATA_BITWIDTH'b11111_11010111000,
        `W_DATA_BITWIDTH'b00000_00101101111,
        `W_DATA_BITWIDTH'b00000_00101011111,
        `W_DATA_BITWIDTH'b11111_11101011010,
        `W_DATA_BITWIDTH'b00000_00100010111,
        `W_DATA_BITWIDTH'b11111_11101110011,
        `W_DATA_BITWIDTH'b11111_11101100010,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b11111_11100110100,
        `W_DATA_BITWIDTH'b11111_11101110000,
        `W_DATA_BITWIDTH'b11111_10111100100,
        `W_DATA_BITWIDTH'b11111_11101011111,
        `W_DATA_BITWIDTH'b00000_00011100101,
        `W_DATA_BITWIDTH'b00000_00100001110,
        `W_DATA_BITWIDTH'b11111_10110010110,
        `W_DATA_BITWIDTH'b00000_00010110000,
        `W_DATA_BITWIDTH'b11111_11101110010,
        `W_DATA_BITWIDTH'b00000_00110001000,
        `W_DATA_BITWIDTH'b11111_11011101011,
        `W_DATA_BITWIDTH'b11111_11101000101,
        `W_DATA_BITWIDTH'b11111_11010001111,
        `W_DATA_BITWIDTH'b00000_00110010101,
        `W_DATA_BITWIDTH'b00000_00010101111,
        `W_DATA_BITWIDTH'b00000_00100000000,
        `W_DATA_BITWIDTH'b11111_11001010000,
        `W_DATA_BITWIDTH'b00000_00011111101,
        `W_DATA_BITWIDTH'b00000_00010101101,
        `W_DATA_BITWIDTH'b00000_00010011100,
        `W_DATA_BITWIDTH'b11111_11101111011,
        `W_DATA_BITWIDTH'b00000_00010110100,
        `W_DATA_BITWIDTH'b11111_11101001010,
        `W_DATA_BITWIDTH'b00000_00011110101,
        `W_DATA_BITWIDTH'b00000_00100111110,
        `W_DATA_BITWIDTH'b00000_00100011011,
        `W_DATA_BITWIDTH'b00000_00010100011,
        `W_DATA_BITWIDTH'b00000_00010001111,
        `W_DATA_BITWIDTH'b11111_11011110101,
        `W_DATA_BITWIDTH'b11111_11100110000,
        `W_DATA_BITWIDTH'b11111_11001100110,
        `W_DATA_BITWIDTH'b00000_00011101101,
        `W_DATA_BITWIDTH'b11111_11100110110,
        `W_DATA_BITWIDTH'b00000_00010110100,
        `W_DATA_BITWIDTH'b11111_11001111101,
        `W_DATA_BITWIDTH'b11111_11011000000,
        `W_DATA_BITWIDTH'b11111_11101010100,
        `W_DATA_BITWIDTH'b11111_11010011000,
        `W_DATA_BITWIDTH'b00000_00011001001,
        `W_DATA_BITWIDTH'b11111_11101010100,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b00000_00010011010,
        `W_DATA_BITWIDTH'b00000_00100010001,
        `W_DATA_BITWIDTH'b11111_11011011011,
        `W_DATA_BITWIDTH'b00000_00010101110,
        `W_DATA_BITWIDTH'b11111_11011011001,
        `W_DATA_BITWIDTH'b00000_00010100011,
        `W_DATA_BITWIDTH'b11111_11101011011,
        `W_DATA_BITWIDTH'b11111_11011000000,
        `W_DATA_BITWIDTH'b11111_11011100111,
        `W_DATA_BITWIDTH'b00000_00011111110,
        `W_DATA_BITWIDTH'b00000_00100000100,
        `W_DATA_BITWIDTH'b00000_00010100100,
        `W_DATA_BITWIDTH'b00000_00011000101,
        `W_DATA_BITWIDTH'b00000_00010000001,
        `W_DATA_BITWIDTH'b00000_00011110100,
        `W_DATA_BITWIDTH'b00000_00010010000,
        `W_DATA_BITWIDTH'b00000_00010111000,
        `W_DATA_BITWIDTH'b00000_00100010000,
        `W_DATA_BITWIDTH'b00000_00100010000,
        `W_DATA_BITWIDTH'b00000_00010001010,
        `W_DATA_BITWIDTH'b00000_00010001101,
        `W_DATA_BITWIDTH'b00000_00010011100,
        `W_DATA_BITWIDTH'b11111_11101100111,
        `W_DATA_BITWIDTH'b11111_10111010111,
        `W_DATA_BITWIDTH'b11111_11001100011,
        `W_DATA_BITWIDTH'b11111_10111111111,
        `W_DATA_BITWIDTH'b11111_10110100011,
        `W_DATA_BITWIDTH'b00000_00010110110,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b00000_00101110000,
        `W_DATA_BITWIDTH'b11111_11010110011,
        `W_DATA_BITWIDTH'b11111_11101100010,
        `W_DATA_BITWIDTH'b11111_10111001110,
        `W_DATA_BITWIDTH'b11111_10001110100,
        `W_DATA_BITWIDTH'b11111_11011001111,
        `W_DATA_BITWIDTH'b00000_00010000010,
        `W_DATA_BITWIDTH'b11111_11101110101,
        `W_DATA_BITWIDTH'b11111_10110011011,
        `W_DATA_BITWIDTH'b11111_11011111001,
        `W_DATA_BITWIDTH'b11111_11011111000,
        `W_DATA_BITWIDTH'b00000_00100011100,
        `W_DATA_BITWIDTH'b11111_11000001101,
        `W_DATA_BITWIDTH'b00000_00100001001,
        `W_DATA_BITWIDTH'b00000_00100111100,
        `W_DATA_BITWIDTH'b00000_00101100110,
        `W_DATA_BITWIDTH'b00000_00101100101,
        `W_DATA_BITWIDTH'b11111_11000010001,
        `W_DATA_BITWIDTH'b00000_00110110101,
        `W_DATA_BITWIDTH'b00000_01000001111,
        `W_DATA_BITWIDTH'b00000_00111011010,
        `W_DATA_BITWIDTH'b11111_11010100100,
        `W_DATA_BITWIDTH'b11111_11100001000,
        `W_DATA_BITWIDTH'b00000_00010001110,
        `W_DATA_BITWIDTH'b11111_11011101111,
        `W_DATA_BITWIDTH'b11111_11011001101,
        `W_DATA_BITWIDTH'b11111_11100010001,
        `W_DATA_BITWIDTH'b00000_00010110000,
        `W_DATA_BITWIDTH'b00000_00101010000,
        `W_DATA_BITWIDTH'b00000_00101010000
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
    '{
        `W_DATA_BITWIDTH'b11111_11101110101,
        `W_DATA_BITWIDTH'b11111_11100100001,
        `W_DATA_BITWIDTH'b11111_11011010011,
        `W_DATA_BITWIDTH'b11111_11010000100,
        `W_DATA_BITWIDTH'b00000_00010100110,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b11111_11011111100,
        `W_DATA_BITWIDTH'b11111_11101100011,
        `W_DATA_BITWIDTH'b11111_11001011101,
        `W_DATA_BITWIDTH'b11111_11100010101,
        `W_DATA_BITWIDTH'b11111_11101010011,
        `W_DATA_BITWIDTH'b11111_11100000110,
        `W_DATA_BITWIDTH'b11111_11001111001,
        `W_DATA_BITWIDTH'b11111_11101100110,
        `W_DATA_BITWIDTH'b00000_00100011111,
        `W_DATA_BITWIDTH'b11111_11010000001,
        `W_DATA_BITWIDTH'b00000_00011111001,
        `W_DATA_BITWIDTH'b11111_11100000010,
        `W_DATA_BITWIDTH'b00000_00010111101,
        `W_DATA_BITWIDTH'b11111_11100100010,
        `W_DATA_BITWIDTH'b00000_00100001111,
        `W_DATA_BITWIDTH'b00000_00010110010,
        `W_DATA_BITWIDTH'b11111_11101100101,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b00000_00011101011,
        `W_DATA_BITWIDTH'b00000_00100100110,
        `W_DATA_BITWIDTH'b00000_00010111100,
        `W_DATA_BITWIDTH'b11111_11101100101,
        `W_DATA_BITWIDTH'b11111_11010111001,
        `W_DATA_BITWIDTH'b11111_11101000101,
        `W_DATA_BITWIDTH'b11111_11100001100,
        `W_DATA_BITWIDTH'b11111_11010011111,
        `W_DATA_BITWIDTH'b00000_00011000111,
        `W_DATA_BITWIDTH'b00000_00011001011,
        `W_DATA_BITWIDTH'b11111_11101010000,
        `W_DATA_BITWIDTH'b00000_00011010100,
        `W_DATA_BITWIDTH'b00000_00010000101,
        `W_DATA_BITWIDTH'b00000_00011111010,
        `W_DATA_BITWIDTH'b11111_11010011010,
        `W_DATA_BITWIDTH'b00000_00010010001,
        `W_DATA_BITWIDTH'b00000_00011010010,
        `W_DATA_BITWIDTH'b00000_00010010100,
        `W_DATA_BITWIDTH'b00000_00010111010,
        `W_DATA_BITWIDTH'b00000_00011111010,
        `W_DATA_BITWIDTH'b11111_11100100011,
        `W_DATA_BITWIDTH'b00000_00010101110,
        `W_DATA_BITWIDTH'b00000_00100111100,
        `W_DATA_BITWIDTH'b11111_11101010101,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b11111_11101000111,
        `W_DATA_BITWIDTH'b00000_00011111010,
        `W_DATA_BITWIDTH'b00000_00011000001,
        `W_DATA_BITWIDTH'b00000_00101000101,
        `W_DATA_BITWIDTH'b11111_11011010000,
        `W_DATA_BITWIDTH'b11111_11001101011,
        `W_DATA_BITWIDTH'b11111_11010100111,
        `W_DATA_BITWIDTH'b11111_11011010001,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b00000_00110101011,
        `W_DATA_BITWIDTH'b00000_00011011010,
        `W_DATA_BITWIDTH'b00000_00100010010,
        `W_DATA_BITWIDTH'b00000_00101000000,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b00000_00100111011,
        `W_DATA_BITWIDTH'b11111_11010110001,
        `W_DATA_BITWIDTH'b11111_11010100001,
        `W_DATA_BITWIDTH'b00000_00101000010,
        `W_DATA_BITWIDTH'b11111_11011101001,
        `W_DATA_BITWIDTH'b11111_11101110101,
        `W_DATA_BITWIDTH'b11111_11010110110,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b00000_00010111011,
        `W_DATA_BITWIDTH'b11111_11010010010,
        `W_DATA_BITWIDTH'b00000_00011111001,
        `W_DATA_BITWIDTH'b00000_00011111001,
        `W_DATA_BITWIDTH'b11111_11001111101,
        `W_DATA_BITWIDTH'b00000_00011101000,
        `W_DATA_BITWIDTH'b11111_11100001110,
        `W_DATA_BITWIDTH'b00000_00101011110,
        `W_DATA_BITWIDTH'b11111_10111101100,
        `W_DATA_BITWIDTH'b00000_00110101001,
        `W_DATA_BITWIDTH'b00000_00011000101,
        `W_DATA_BITWIDTH'b00000_00100110111,
        `W_DATA_BITWIDTH'b11111_10100110000,
        `W_DATA_BITWIDTH'b00000_00110000111,
        `W_DATA_BITWIDTH'b11111_11011100010,
        `W_DATA_BITWIDTH'b11111_11010000110,
        `W_DATA_BITWIDTH'b11111_11001000001,
        `W_DATA_BITWIDTH'b11111_10100100101,
        `W_DATA_BITWIDTH'b11111_11100101100,
        `W_DATA_BITWIDTH'b11111_11001000111,
        `W_DATA_BITWIDTH'b00000_00011010110,
        `W_DATA_BITWIDTH'b00000_00110101010,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b11111_11100000111,
        `W_DATA_BITWIDTH'b11111_11100111011,
        `W_DATA_BITWIDTH'b11111_11000001100,
        `W_DATA_BITWIDTH'b00000_00101100111,
        `W_DATA_BITWIDTH'b00000_00111111010,
        `W_DATA_BITWIDTH'b00000_00111010110,
        `W_DATA_BITWIDTH'b00000_00010110100,
        `W_DATA_BITWIDTH'b00000_00101001011,
        `W_DATA_BITWIDTH'b00000_00111111000,
        `W_DATA_BITWIDTH'b00000_00010111101,
        `W_DATA_BITWIDTH'b00000_00101001000,
        `W_DATA_BITWIDTH'b11111_10100110011,
        `W_DATA_BITWIDTH'b00000_00110100100,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b11111_11011001001,
        `W_DATA_BITWIDTH'b00000_01001110111,
        `W_DATA_BITWIDTH'b00000_01001011010,
        `W_DATA_BITWIDTH'b00000_00011001001,
        `W_DATA_BITWIDTH'b11111_11011101100,
        `W_DATA_BITWIDTH'b11111_11001110110,
        `W_DATA_BITWIDTH'b00000_00010000101,
        `W_DATA_BITWIDTH'b11111_11000101001,
        `W_DATA_BITWIDTH'b11111_11001100101,
        `W_DATA_BITWIDTH'b00000_00101101010,
        `W_DATA_BITWIDTH'b11111_11100111010,
        `W_DATA_BITWIDTH'b11111_11001001101,
        `W_DATA_BITWIDTH'b11111_11101011101,
        `W_DATA_BITWIDTH'b00000_00011010111,
        `W_DATA_BITWIDTH'b11111_10111000101,
        `W_DATA_BITWIDTH'b00000_00010101110,
        `W_DATA_BITWIDTH'b00000_00100000101,
        `W_DATA_BITWIDTH'b11111_11101111111,
        `W_DATA_BITWIDTH'b11111_11100111001,
        `W_DATA_BITWIDTH'b11111_11011100011,
        `W_DATA_BITWIDTH'b11111_11101001001,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b00000_00011010010,
        `W_DATA_BITWIDTH'b11111_11100100100,
        `W_DATA_BITWIDTH'b11111_11011110000,
        `W_DATA_BITWIDTH'b11111_11011110011,
        `W_DATA_BITWIDTH'b11111_11101111010,
        `W_DATA_BITWIDTH'b00000_00011110010,
        `W_DATA_BITWIDTH'b00000_00010100011,
        `W_DATA_BITWIDTH'b11111_11000110011,
        `W_DATA_BITWIDTH'b00000_00101110101,
        `W_DATA_BITWIDTH'b00000_00010100111,
        `W_DATA_BITWIDTH'b11111_11101010000,
        `W_DATA_BITWIDTH'b00000_00100001111,
        `W_DATA_BITWIDTH'b00000_00010101001,
        `W_DATA_BITWIDTH'b00000_00010101011,
        `W_DATA_BITWIDTH'b11111_11100110111,
        `W_DATA_BITWIDTH'b00000_00011000111,
        `W_DATA_BITWIDTH'b11111_11011110001,
        `W_DATA_BITWIDTH'b00000_00100100110,
        `W_DATA_BITWIDTH'b11111_11000010011,
        `W_DATA_BITWIDTH'b11111_11100001001,
        `W_DATA_BITWIDTH'b11111_11101000001,
        `W_DATA_BITWIDTH'b11111_11100011111,
        `W_DATA_BITWIDTH'b11111_11100101011,
        `W_DATA_BITWIDTH'b11111_11101101101,
        `W_DATA_BITWIDTH'b11111_11100011010,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b00000_00100110011,
        `W_DATA_BITWIDTH'b00000_00100010110,
        `W_DATA_BITWIDTH'b00000_00010000001,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b11111_11100010001,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b00000_00011101110,
        `W_DATA_BITWIDTH'b11111_11100110101,
        `W_DATA_BITWIDTH'b00000_00010101001,
        `W_DATA_BITWIDTH'b00000_00011101011,
        `W_DATA_BITWIDTH'b00000_00010011111,
        `W_DATA_BITWIDTH'b11111_11011000010,
        `W_DATA_BITWIDTH'b00000_00010010101,
        `W_DATA_BITWIDTH'b00000_00011001000,
        `W_DATA_BITWIDTH'b00000_00010001000,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b00000_00010101101,
        `W_DATA_BITWIDTH'b11111_11011100100,
        `W_DATA_BITWIDTH'b00000_00011001010,
        `W_DATA_BITWIDTH'b11111_11101001001,
        `W_DATA_BITWIDTH'b00000_00011010011,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b11111_11100001000,
        `W_DATA_BITWIDTH'b11111_11011010111,
        `W_DATA_BITWIDTH'b00000_00011100001,
        `W_DATA_BITWIDTH'b00000_00101110111,
        `W_DATA_BITWIDTH'b00000_00010100111,
        `W_DATA_BITWIDTH'b00000_00010001100,
        `W_DATA_BITWIDTH'b11111_11011010101,
        `W_DATA_BITWIDTH'b11111_11101111010,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b00000_00010000101,
        `W_DATA_BITWIDTH'b00000_00101110001,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b00000_00100001110,
        `W_DATA_BITWIDTH'b11111_11011000010,
        `W_DATA_BITWIDTH'b11111_11011100100,
        `W_DATA_BITWIDTH'b11111_11101110100,
        `W_DATA_BITWIDTH'b11111_11101101110,
        `W_DATA_BITWIDTH'b11111_11101001000,
        `W_DATA_BITWIDTH'b00000_00010101110,
        `W_DATA_BITWIDTH'b11111_11101010010,
        `W_DATA_BITWIDTH'b11111_11001110010,
        `W_DATA_BITWIDTH'b00000_00010100000,
        `W_DATA_BITWIDTH'b11111_11100011100,
        `W_DATA_BITWIDTH'b00000_00011110110,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b00000_00011001100,
        `W_DATA_BITWIDTH'b11111_11101011011,
        `W_DATA_BITWIDTH'b00000_00010101001,
        `W_DATA_BITWIDTH'b11111_11100010110,
        `W_DATA_BITWIDTH'b11111_11011110001,
        `W_DATA_BITWIDTH'b11111_11001010000,
        `W_DATA_BITWIDTH'b11111_11011111111,
        `W_DATA_BITWIDTH'b00000_00011001000,
        `W_DATA_BITWIDTH'b11111_11011100011,
        `W_DATA_BITWIDTH'b11111_11100111000,
        `W_DATA_BITWIDTH'b11111_11100110100,
        `W_DATA_BITWIDTH'b11111_11010110010,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b00000_00011101001,
        `W_DATA_BITWIDTH'b11111_11100010111,
        `W_DATA_BITWIDTH'b11111_11101110111,
        `W_DATA_BITWIDTH'b00000_00011010010,
        `W_DATA_BITWIDTH'b00000_00110010010,
        `W_DATA_BITWIDTH'b00000_00011110101,
        `W_DATA_BITWIDTH'b11111_11101010110,
        `W_DATA_BITWIDTH'b00000_00010101000,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b00000_00100000100,
        `W_DATA_BITWIDTH'b00000_00011000011,
        `W_DATA_BITWIDTH'b00000_00111101000,
        `W_DATA_BITWIDTH'b00000_01000111011,
        `W_DATA_BITWIDTH'b00000_00111010000,
        `W_DATA_BITWIDTH'b00000_00010111111,
        `W_DATA_BITWIDTH'b11111_11101100000,
        `W_DATA_BITWIDTH'b00000_00101100011,
        `W_DATA_BITWIDTH'b11111_10110110001,
        `W_DATA_BITWIDTH'b00000_01000011111,
        `W_DATA_BITWIDTH'b11111_11100101011,
        `W_DATA_BITWIDTH'b11111_11000011100,
        `W_DATA_BITWIDTH'b00000_00111110101,
        `W_DATA_BITWIDTH'b11111_11100110000,
        `W_DATA_BITWIDTH'b11111_11010111000,
        `W_DATA_BITWIDTH'b11111_10110101110,
        `W_DATA_BITWIDTH'b00000_00101000001,
        `W_DATA_BITWIDTH'b00000_00110100011,
        `W_DATA_BITWIDTH'b00000_00100111011,
        `W_DATA_BITWIDTH'b00000_00100001000,
        `W_DATA_BITWIDTH'b11111_10101001010,
        `W_DATA_BITWIDTH'b11111_11000101010,
        `W_DATA_BITWIDTH'b00000_00101001100,
        `W_DATA_BITWIDTH'b00000_00100000101,
        `W_DATA_BITWIDTH'b11111_11100110000,
        `W_DATA_BITWIDTH'b00000_00011100100,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b11111_10111010001,
        `W_DATA_BITWIDTH'b11111_11101000111,
        `W_DATA_BITWIDTH'b00000_00011110100,
        `W_DATA_BITWIDTH'b00000_00110101110,
        `W_DATA_BITWIDTH'b11111_11100110110,
        `W_DATA_BITWIDTH'b00000_00100100111,
        `W_DATA_BITWIDTH'b11111_10111010011,
        `W_DATA_BITWIDTH'b00000_00110101101,
        `W_DATA_BITWIDTH'b00000_00011010110,
        `W_DATA_BITWIDTH'b00000_00101110110,
        `W_DATA_BITWIDTH'b11111_11101011010,
        `W_DATA_BITWIDTH'b00000_00010011000,
        `W_DATA_BITWIDTH'b00000_00011100000,
        `W_DATA_BITWIDTH'b11111_11100111110,
        `W_DATA_BITWIDTH'b11111_11100011101,
        `W_DATA_BITWIDTH'b11111_11101101111,
        `W_DATA_BITWIDTH'b00000_00010111111,
        `W_DATA_BITWIDTH'b00000_00011011101,
        `W_DATA_BITWIDTH'b11111_11100000011,
        `W_DATA_BITWIDTH'b11111_11011101111,
        `W_DATA_BITWIDTH'b00000_00011011101,
        `W_DATA_BITWIDTH'b00000_00010110100,
        `W_DATA_BITWIDTH'b11111_11101010010,
        `W_DATA_BITWIDTH'b11111_11010010101,
        `W_DATA_BITWIDTH'b00000_00100001111,
        `W_DATA_BITWIDTH'b00000_00100111010,
        `W_DATA_BITWIDTH'b00000_00010110001,
        `W_DATA_BITWIDTH'b00000_00010000110,
        `W_DATA_BITWIDTH'b00000_00010101111,
        `W_DATA_BITWIDTH'b00000_00110111111,
        `W_DATA_BITWIDTH'b11111_11100000000,
        `W_DATA_BITWIDTH'b11111_11101100000,
        `W_DATA_BITWIDTH'b11111_11100011101,
        `W_DATA_BITWIDTH'b00000_01000011001,
        `W_DATA_BITWIDTH'b11111_11010001010,
        `W_DATA_BITWIDTH'b11111_11011001111,
        `W_DATA_BITWIDTH'b11111_11100101100,
        `W_DATA_BITWIDTH'b11111_11001110110,
        `W_DATA_BITWIDTH'b00000_00011111101,
        `W_DATA_BITWIDTH'b00000_00100110101,
        `W_DATA_BITWIDTH'b11111_11000111011,
        `W_DATA_BITWIDTH'b00000_00010000001,
        `W_DATA_BITWIDTH'b00000_00011010110,
        `W_DATA_BITWIDTH'b11111_11011101111,
        `W_DATA_BITWIDTH'b00000_00010000010,
        `W_DATA_BITWIDTH'b11111_11010010011,
        `W_DATA_BITWIDTH'b11111_11100111010,
        `W_DATA_BITWIDTH'b11111_11011111110,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b11111_11100001001,
        `W_DATA_BITWIDTH'b00000_00010011000,
        `W_DATA_BITWIDTH'b00000_00010011010,
        `W_DATA_BITWIDTH'b11111_11100101101,
        `W_DATA_BITWIDTH'b00000_00011100100,
        `W_DATA_BITWIDTH'b11111_11001110100,
        `W_DATA_BITWIDTH'b11111_11001001011,
        `W_DATA_BITWIDTH'b00000_00100110101,
        `W_DATA_BITWIDTH'b11111_11011010100,
        `W_DATA_BITWIDTH'b00000_01000110110,
        `W_DATA_BITWIDTH'b00000_00101100111,
        `W_DATA_BITWIDTH'b00000_00101010011,
        `W_DATA_BITWIDTH'b11111_11001110111,
        `W_DATA_BITWIDTH'b11111_11101000001,
        `W_DATA_BITWIDTH'b00000_00101111101,
        `W_DATA_BITWIDTH'b11111_11010000100,
        `W_DATA_BITWIDTH'b00000_00110011110,
        `W_DATA_BITWIDTH'b00000_00101010101,
        `W_DATA_BITWIDTH'b00000_00100100000,
        `W_DATA_BITWIDTH'b11111_11010100000,
        `W_DATA_BITWIDTH'b11111_10110011101,
        `W_DATA_BITWIDTH'b11111_11101000001,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b00000_00010110100,
        `W_DATA_BITWIDTH'b11111_11100000101,
        `W_DATA_BITWIDTH'b11111_10010111001,
        `W_DATA_BITWIDTH'b00000_01000011100,
        `W_DATA_BITWIDTH'b00000_00010110110,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b11111_11100010000,
        `W_DATA_BITWIDTH'b11111_10010011011,
        `W_DATA_BITWIDTH'b00000_00010000110,
        `W_DATA_BITWIDTH'b11111_10101111011,
        `W_DATA_BITWIDTH'b11111_11001101010,
        `W_DATA_BITWIDTH'b00000_00111010110,
        `W_DATA_BITWIDTH'b11111_11100100001,
        `W_DATA_BITWIDTH'b11111_11000100001,
        `W_DATA_BITWIDTH'b11111_11001011001,
        `W_DATA_BITWIDTH'b11111_11010111100,
        `W_DATA_BITWIDTH'b11111_11000101001,
        `W_DATA_BITWIDTH'b00000_00010001111,
        `W_DATA_BITWIDTH'b11111_11001000101,
        `W_DATA_BITWIDTH'b00000_00010010010,
        `W_DATA_BITWIDTH'b11111_11011000000,
        `W_DATA_BITWIDTH'b00000_00010011111,
        `W_DATA_BITWIDTH'b11111_11101001000,
        `W_DATA_BITWIDTH'b11111_11101101010,
        `W_DATA_BITWIDTH'b00000_00010011110,
        `W_DATA_BITWIDTH'b11111_11011000001,
        `W_DATA_BITWIDTH'b11111_11010110011,
        `W_DATA_BITWIDTH'b11111_11101100011,
        `W_DATA_BITWIDTH'b00000_00100011011,
        `W_DATA_BITWIDTH'b11111_11000110110,
        `W_DATA_BITWIDTH'b11111_11101100011,
        `W_DATA_BITWIDTH'b11111_11000010011,
        `W_DATA_BITWIDTH'b11111_11100100101,
        `W_DATA_BITWIDTH'b11111_11100101101,
        `W_DATA_BITWIDTH'b00000_00110010110,
        `W_DATA_BITWIDTH'b00000_00010110101,
        `W_DATA_BITWIDTH'b11111_11101001011,
        `W_DATA_BITWIDTH'b11111_11101010100,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b00000_00011001000,
        `W_DATA_BITWIDTH'b11111_11101100100,
        `W_DATA_BITWIDTH'b00000_00010100001,
        `W_DATA_BITWIDTH'b00000_00010000110,
        `W_DATA_BITWIDTH'b11111_11100101110,
        `W_DATA_BITWIDTH'b11111_11100111111,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b11111_11001100011,
        `W_DATA_BITWIDTH'b00000_00110011110,
        `W_DATA_BITWIDTH'b00000_00101110111,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b00000_00011000011,
        `W_DATA_BITWIDTH'b11111_11101101111,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b00000_00100101111,
        `W_DATA_BITWIDTH'b11111_11101100001,
        `W_DATA_BITWIDTH'b00000_00101110000,
        `W_DATA_BITWIDTH'b00000_00101010010,
        `W_DATA_BITWIDTH'b00000_00110000111,
        `W_DATA_BITWIDTH'b00000_00011000101,
        `W_DATA_BITWIDTH'b00000_00100111110,
        `W_DATA_BITWIDTH'b00000_00010001011,
        `W_DATA_BITWIDTH'b11111_11010110101,
        `W_DATA_BITWIDTH'b11111_11101111011,
        `W_DATA_BITWIDTH'b00000_00100010101,
        `W_DATA_BITWIDTH'b11111_11011001111,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b00000_00100001011,
        `W_DATA_BITWIDTH'b00000_00010001001,
        `W_DATA_BITWIDTH'b11111_11100100000,
        `W_DATA_BITWIDTH'b00000_00100000001,
        `W_DATA_BITWIDTH'b00000_00100111111,
        `W_DATA_BITWIDTH'b11111_11010101010,
        `W_DATA_BITWIDTH'b00000_00010110001,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b11111_10110110000,
        `W_DATA_BITWIDTH'b11111_11101000011,
        `W_DATA_BITWIDTH'b11111_11101110111,
        `W_DATA_BITWIDTH'b00000_00011001100,
        `W_DATA_BITWIDTH'b00000_00010101010,
        `W_DATA_BITWIDTH'b00000_00010001100,
        `W_DATA_BITWIDTH'b11111_11101110111,
        `W_DATA_BITWIDTH'b11111_11011110001,
        `W_DATA_BITWIDTH'b00000_00011001101,
        `W_DATA_BITWIDTH'b00000_00100100110,
        `W_DATA_BITWIDTH'b11111_11101110000,
        `W_DATA_BITWIDTH'b11111_11100110010,
        `W_DATA_BITWIDTH'b00000_00010010101,
        `W_DATA_BITWIDTH'b00000_00101010110,
        `W_DATA_BITWIDTH'b00000_00011011000,
        `W_DATA_BITWIDTH'b00000_00010111101,
        `W_DATA_BITWIDTH'b00000_00010110100,
        `W_DATA_BITWIDTH'b00000_00011100010,
        `W_DATA_BITWIDTH'b11111_11101110100,
        `W_DATA_BITWIDTH'b00000_00010101101,
        `W_DATA_BITWIDTH'b00000_00010000100,
        `W_DATA_BITWIDTH'b00000_00010111010,
        `W_DATA_BITWIDTH'b00000_00100100010,
        `W_DATA_BITWIDTH'b00000_00011010111,
        `W_DATA_BITWIDTH'b00000_00010111011,
        `W_DATA_BITWIDTH'b00000_00100000101,
        `W_DATA_BITWIDTH'b11111_11100000101,
        `W_DATA_BITWIDTH'b11111_10110010000,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b11111_11011111011,
        `W_DATA_BITWIDTH'b11111_11011100001,
        `W_DATA_BITWIDTH'b00000_00101011000,
        `W_DATA_BITWIDTH'b00000_00010000001,
        `W_DATA_BITWIDTH'b00000_00011011000,
        `W_DATA_BITWIDTH'b11111_11101110101,
        `W_DATA_BITWIDTH'b11111_10110101100,
        `W_DATA_BITWIDTH'b11111_11100010110,
        `W_DATA_BITWIDTH'b11111_11100001100,
        `W_DATA_BITWIDTH'b11111_11100100101,
        `W_DATA_BITWIDTH'b11111_11100011011,
        `W_DATA_BITWIDTH'b00000_00010111010,
        `W_DATA_BITWIDTH'b11111_11010001110,
        `W_DATA_BITWIDTH'b11111_11100001110,
        `W_DATA_BITWIDTH'b00000_00011101011,
        `W_DATA_BITWIDTH'b11111_11000010010,
        `W_DATA_BITWIDTH'b00000_00100010111,
        `W_DATA_BITWIDTH'b11111_11010001110,
        `W_DATA_BITWIDTH'b11111_11010110101,
        `W_DATA_BITWIDTH'b00000_00010111111,
        `W_DATA_BITWIDTH'b00000_00010001111,
        `W_DATA_BITWIDTH'b11111_11100000101,
        `W_DATA_BITWIDTH'b11111_11000000110,
        `W_DATA_BITWIDTH'b11111_11101100010,
        `W_DATA_BITWIDTH'b11111_11010100100,
        `W_DATA_BITWIDTH'b00000_00100100010,
        `W_DATA_BITWIDTH'b00000_00110000001,
        `W_DATA_BITWIDTH'b00000_00100000000,
        `W_DATA_BITWIDTH'b00000_01001000010,
        `W_DATA_BITWIDTH'b00000_01001000010
    };
    localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
    '{
        `W_DATA_BITWIDTH'b00000_00010100010,
        `W_DATA_BITWIDTH'b11111_11100010000,
        `W_DATA_BITWIDTH'b00000_00011010101,
        `W_DATA_BITWIDTH'b11111_11011000000,
        `W_DATA_BITWIDTH'b11111_11101100100,
        `W_DATA_BITWIDTH'b00000_00011010001,
        `W_DATA_BITWIDTH'b00000_00011110111,
        `W_DATA_BITWIDTH'b00000_00011010100,
        `W_DATA_BITWIDTH'b11111_11011110100,
        `W_DATA_BITWIDTH'b11111_11010010100,
        `W_DATA_BITWIDTH'b00000_00010010010,
        `W_DATA_BITWIDTH'b11111_11001110100,
        `W_DATA_BITWIDTH'b00000_00011111100,
        `W_DATA_BITWIDTH'b00000_00011000111,
        `W_DATA_BITWIDTH'b11111_11100111010,
        `W_DATA_BITWIDTH'b11111_11101110111,
        `W_DATA_BITWIDTH'b00000_00010011000,
        `W_DATA_BITWIDTH'b11111_11100011011,
        `W_DATA_BITWIDTH'b00000_00100110101,
        `W_DATA_BITWIDTH'b11111_11011111001,
        `W_DATA_BITWIDTH'b11111_11100000010,
        `W_DATA_BITWIDTH'b00000_00101001111,
        `W_DATA_BITWIDTH'b11111_11101011000,
        `W_DATA_BITWIDTH'b00000_00100000010,
        `W_DATA_BITWIDTH'b11111_11100101010,
        `W_DATA_BITWIDTH'b11111_11011001011,
        `W_DATA_BITWIDTH'b11111_11100100110,
        `W_DATA_BITWIDTH'b00000_00010010000,
        `W_DATA_BITWIDTH'b00000_00010000100,
        `W_DATA_BITWIDTH'b11111_11011111100,
        `W_DATA_BITWIDTH'b11111_11010110001,
        `W_DATA_BITWIDTH'b11111_11011001111,
        `W_DATA_BITWIDTH'b11111_11101110101,
        `W_DATA_BITWIDTH'b00000_00100101100,
        `W_DATA_BITWIDTH'b00000_00010101010,
        `W_DATA_BITWIDTH'b00000_00100101011,
        `W_DATA_BITWIDTH'b11111_11101010011,
        `W_DATA_BITWIDTH'b11111_11101100011,
        `W_DATA_BITWIDTH'b11111_11100000000,
        `W_DATA_BITWIDTH'b11111_11010110010,
        `W_DATA_BITWIDTH'b11111_11010000100,
        `W_DATA_BITWIDTH'b11111_11101000110,
        `W_DATA_BITWIDTH'b00000_00010101000,
        `W_DATA_BITWIDTH'b00000_00010010111,
        `W_DATA_BITWIDTH'b00000_00101000111,
        `W_DATA_BITWIDTH'b00000_01000110101,
        `W_DATA_BITWIDTH'b11111_11010010101,
        `W_DATA_BITWIDTH'b00000_00010010110,
        `W_DATA_BITWIDTH'b00000_00011111111,
        `W_DATA_BITWIDTH'b00000_00011100110,
        `W_DATA_BITWIDTH'b11111_11010000101,
        `W_DATA_BITWIDTH'b00000_00010101100,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b00000_00010001101,
        `W_DATA_BITWIDTH'b00000_00011101010,
        `W_DATA_BITWIDTH'b11111_11101110001,
        `W_DATA_BITWIDTH'b00000_00011100111,
        `W_DATA_BITWIDTH'b11111_11101011010,
        `W_DATA_BITWIDTH'b00000_00011011010,
        `W_DATA_BITWIDTH'b11111_11100111011,
        `W_DATA_BITWIDTH'b11111_11101110010,
        `W_DATA_BITWIDTH'b11111_11100111111,
        `W_DATA_BITWIDTH'b00000_00100010000,
        `W_DATA_BITWIDTH'b11111_11100111000,
        `W_DATA_BITWIDTH'b00000_00011111100,
        `W_DATA_BITWIDTH'b00000_00011101100,
        `W_DATA_BITWIDTH'b00000_00100011001,
        `W_DATA_BITWIDTH'b11111_11000101110,
        `W_DATA_BITWIDTH'b00000_00111111110,
        `W_DATA_BITWIDTH'b11111_11001111000,
        `W_DATA_BITWIDTH'b11111_11100110011,
        `W_DATA_BITWIDTH'b11111_11000101101,
        `W_DATA_BITWIDTH'b00000_00011000011,
        `W_DATA_BITWIDTH'b11111_10111100011,
        `W_DATA_BITWIDTH'b11111_11011001111,
        `W_DATA_BITWIDTH'b00000_01011111010,
        `W_DATA_BITWIDTH'b00000_00100011000,
        `W_DATA_BITWIDTH'b00000_00110000001,
        `W_DATA_BITWIDTH'b11111_11011100101,
        `W_DATA_BITWIDTH'b11111_11010110001,
        `W_DATA_BITWIDTH'b00000_00010101011,
        `W_DATA_BITWIDTH'b11111_10111100100,
        `W_DATA_BITWIDTH'b11111_11101111010,
        `W_DATA_BITWIDTH'b11111_11101111001,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b00000_00010011111,
        `W_DATA_BITWIDTH'b00000_00101101110,
        `W_DATA_BITWIDTH'b00000_00011111110,
        `W_DATA_BITWIDTH'b00000_01000101110,
        `W_DATA_BITWIDTH'b11111_11000011001,
        `W_DATA_BITWIDTH'b00000_00100000001,
        `W_DATA_BITWIDTH'b00000_00101010111,
        `W_DATA_BITWIDTH'b11111_11001001100,
        `W_DATA_BITWIDTH'b11111_11011111101,
        `W_DATA_BITWIDTH'b11111_11100010001,
        `W_DATA_BITWIDTH'b00000_00110101010,
        `W_DATA_BITWIDTH'b11111_11100111111,
        `W_DATA_BITWIDTH'b11111_11001011101,
        `W_DATA_BITWIDTH'b11111_11100001100,
        `W_DATA_BITWIDTH'b00000_00010101010,
        `W_DATA_BITWIDTH'b11111_10110110001,
        `W_DATA_BITWIDTH'b11111_11101101101,
        `W_DATA_BITWIDTH'b11111_10110111000,
        `W_DATA_BITWIDTH'b00000_01010000111,
        `W_DATA_BITWIDTH'b00000_00010001111,
        `W_DATA_BITWIDTH'b00000_00100100111,
        `W_DATA_BITWIDTH'b00000_00100000001,
        `W_DATA_BITWIDTH'b11111_10110111110,
        `W_DATA_BITWIDTH'b00000_00110101001,
        `W_DATA_BITWIDTH'b11111_11001101010,
        `W_DATA_BITWIDTH'b11111_10100100011,
        `W_DATA_BITWIDTH'b00000_00011101100,
        `W_DATA_BITWIDTH'b11111_11000000111,
        `W_DATA_BITWIDTH'b11111_11100001011,
        `W_DATA_BITWIDTH'b11111_11011010000,
        `W_DATA_BITWIDTH'b11111_11001000101,
        `W_DATA_BITWIDTH'b11111_11101011111,
        `W_DATA_BITWIDTH'b11111_10110100000,
        `W_DATA_BITWIDTH'b11111_11001111111,
        `W_DATA_BITWIDTH'b00000_00101101110,
        `W_DATA_BITWIDTH'b11111_11100100111,
        `W_DATA_BITWIDTH'b11111_11001111010,
        `W_DATA_BITWIDTH'b00000_00010100111,
        `W_DATA_BITWIDTH'b00000_00100010011,
        `W_DATA_BITWIDTH'b11111_11011010001,
        `W_DATA_BITWIDTH'b00000_00101010111,
        `W_DATA_BITWIDTH'b11111_11010111000,
        `W_DATA_BITWIDTH'b11111_11101010111,
        `W_DATA_BITWIDTH'b11111_11100101000,
        `W_DATA_BITWIDTH'b11111_11100010111,
        `W_DATA_BITWIDTH'b00000_00010000010,
        `W_DATA_BITWIDTH'b11111_11100100011,
        `W_DATA_BITWIDTH'b00000_00010011011,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b11111_11100111101,
        `W_DATA_BITWIDTH'b00000_00011000101,
        `W_DATA_BITWIDTH'b00000_00010010111,
        `W_DATA_BITWIDTH'b11111_11101101000,
        `W_DATA_BITWIDTH'b00000_00011111111,
        `W_DATA_BITWIDTH'b00000_00101011001,
        `W_DATA_BITWIDTH'b00000_00011010100,
        `W_DATA_BITWIDTH'b11111_11011110101,
        `W_DATA_BITWIDTH'b11111_11101011001,
        `W_DATA_BITWIDTH'b00000_00010011000,
        `W_DATA_BITWIDTH'b11111_11010001001,
        `W_DATA_BITWIDTH'b00000_00100000111,
        `W_DATA_BITWIDTH'b11111_11101110010,
        `W_DATA_BITWIDTH'b00000_00010011001,
        `W_DATA_BITWIDTH'b11111_11100010011,
        `W_DATA_BITWIDTH'b11111_11001111111,
        `W_DATA_BITWIDTH'b00000_00010100011,
        `W_DATA_BITWIDTH'b11111_11011100000,
        `W_DATA_BITWIDTH'b00000_00101111010,
        `W_DATA_BITWIDTH'b11111_11100101111,
        `W_DATA_BITWIDTH'b11111_11001111010,
        `W_DATA_BITWIDTH'b00000_00011101100,
        `W_DATA_BITWIDTH'b11111_11011001000,
        `W_DATA_BITWIDTH'b11111_11100100000,
        `W_DATA_BITWIDTH'b00000_00011000101,
        `W_DATA_BITWIDTH'b11111_11100001110,
        `W_DATA_BITWIDTH'b00000_00011001000,
        `W_DATA_BITWIDTH'b11111_11001100100,
        `W_DATA_BITWIDTH'b00000_00100100000,
        `W_DATA_BITWIDTH'b11111_11101010000,
        `W_DATA_BITWIDTH'b11111_11001001011,
        `W_DATA_BITWIDTH'b11111_11011110010,
        `W_DATA_BITWIDTH'b11111_10111010100,
        `W_DATA_BITWIDTH'b11111_11011101101,
        `W_DATA_BITWIDTH'b11111_11011001010,
        `W_DATA_BITWIDTH'b11111_11001101101,
        `W_DATA_BITWIDTH'b11111_11101110010,
        `W_DATA_BITWIDTH'b11111_11100010000,
        `W_DATA_BITWIDTH'b00000_00010000100,
        `W_DATA_BITWIDTH'b11111_11100010001,
        `W_DATA_BITWIDTH'b00000_00010011101,
        `W_DATA_BITWIDTH'b00000_00100000101,
        `W_DATA_BITWIDTH'b11111_11100001110,
        `W_DATA_BITWIDTH'b00000_00100111000,
        `W_DATA_BITWIDTH'b11111_11001111100,
        `W_DATA_BITWIDTH'b11111_11101010011,
        `W_DATA_BITWIDTH'b11111_11100101000,
        `W_DATA_BITWIDTH'b11111_11100010001,
        `W_DATA_BITWIDTH'b00000_00011011111,
        `W_DATA_BITWIDTH'b11111_11101010111,
        `W_DATA_BITWIDTH'b11111_11101011010,
        `W_DATA_BITWIDTH'b11111_10111101111,
        `W_DATA_BITWIDTH'b11111_11100111111,
        `W_DATA_BITWIDTH'b11111_11100111101,
        `W_DATA_BITWIDTH'b00000_00010100001,
        `W_DATA_BITWIDTH'b00000_00100100011,
        `W_DATA_BITWIDTH'b00000_00010010011,
        `W_DATA_BITWIDTH'b11111_10110101010,
        `W_DATA_BITWIDTH'b11111_11010011000,
        `W_DATA_BITWIDTH'b00000_00010000100,
        `W_DATA_BITWIDTH'b00000_00101001100,
        `W_DATA_BITWIDTH'b11111_11100100111,
        `W_DATA_BITWIDTH'b11111_11100001010,
        `W_DATA_BITWIDTH'b11111_11001111101,
        `W_DATA_BITWIDTH'b11111_11011011101,
        `W_DATA_BITWIDTH'b11111_11010101100,
        `W_DATA_BITWIDTH'b00000_00010001000,
        `W_DATA_BITWIDTH'b11111_11000110010,
        `W_DATA_BITWIDTH'b00000_00101001100,
        `W_DATA_BITWIDTH'b11111_11011110101,
        `W_DATA_BITWIDTH'b00000_00010000011,
        `W_DATA_BITWIDTH'b00000_00100111010,
        `W_DATA_BITWIDTH'b11111_11011001001,
        `W_DATA_BITWIDTH'b00000_00011111000,
        `W_DATA_BITWIDTH'b00000_00010010111,
        `W_DATA_BITWIDTH'b11111_11011011011,
        `W_DATA_BITWIDTH'b11111_11011000010,
        `W_DATA_BITWIDTH'b11111_11010111111,
        `W_DATA_BITWIDTH'b11111_11011101100,
        `W_DATA_BITWIDTH'b00000_00010001111,
        `W_DATA_BITWIDTH'b11111_11010011101,
        `W_DATA_BITWIDTH'b11111_11101111101,
        `W_DATA_BITWIDTH'b00000_00011101110,
        `W_DATA_BITWIDTH'b00000_00010001011,
        `W_DATA_BITWIDTH'b11111_11100011000,
        `W_DATA_BITWIDTH'b00000_00011000001,
        `W_DATA_BITWIDTH'b11111_11101101000,
        `W_DATA_BITWIDTH'b11111_11101001110,
        `W_DATA_BITWIDTH'b11111_11010110011,
        `W_DATA_BITWIDTH'b00000_00101001100,
        `W_DATA_BITWIDTH'b11111_11010101000,
        `W_DATA_BITWIDTH'b11111_11011110011,
        `W_DATA_BITWIDTH'b11111_11000011101,
        `W_DATA_BITWIDTH'b00000_00010001101,
        `W_DATA_BITWIDTH'b11111_11010100100,
        `W_DATA_BITWIDTH'b00000_00010000010,
        `W_DATA_BITWIDTH'b00000_00010100110,
        `W_DATA_BITWIDTH'b11111_11100111000,
        `W_DATA_BITWIDTH'b00000_00101100101,
        `W_DATA_BITWIDTH'b00000_00101000110,
        `W_DATA_BITWIDTH'b11111_11011011100,
        `W_DATA_BITWIDTH'b00000_00010011111,
        `W_DATA_BITWIDTH'b11111_11000110101,
        `W_DATA_BITWIDTH'b00000_00100100111,
        `W_DATA_BITWIDTH'b11111_10010101100,
        `W_DATA_BITWIDTH'b11111_10101111001,
        `W_DATA_BITWIDTH'b00000_00011100100,
        `W_DATA_BITWIDTH'b11111_11010010111,
        `W_DATA_BITWIDTH'b11111_11001100101,
        `W_DATA_BITWIDTH'b00000_00101010110,
        `W_DATA_BITWIDTH'b00000_00010011001,
        `W_DATA_BITWIDTH'b00000_01010001010,
        `W_DATA_BITWIDTH'b11111_11000111101,
        `W_DATA_BITWIDTH'b00000_00011110011,
        `W_DATA_BITWIDTH'b11111_11001000111,
        `W_DATA_BITWIDTH'b11111_11010100111,
        `W_DATA_BITWIDTH'b11111_11000110000,
        `W_DATA_BITWIDTH'b11111_11000101011,
        `W_DATA_BITWIDTH'b00000_00100100000,
        `W_DATA_BITWIDTH'b00000_00011011011,
        `W_DATA_BITWIDTH'b11111_11100111011,
        `W_DATA_BITWIDTH'b00000_00010001011,
        `W_DATA_BITWIDTH'b00000_00111001010,
        `W_DATA_BITWIDTH'b00000_00101001000,
        `W_DATA_BITWIDTH'b11111_11001011001,
        `W_DATA_BITWIDTH'b00000_00101011010,
        `W_DATA_BITWIDTH'b00000_00011101001,
        `W_DATA_BITWIDTH'b11111_11101111110,
        `W_DATA_BITWIDTH'b11111_11010101010,
        `W_DATA_BITWIDTH'b00000_00011110000,
        `W_DATA_BITWIDTH'b11111_11100101011,
        `W_DATA_BITWIDTH'b00000_00010100110,
        `W_DATA_BITWIDTH'b11111_11100111101,
        `W_DATA_BITWIDTH'b00000_00100001100,
        `W_DATA_BITWIDTH'b00000_00101000100,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b00000_00011001010,
        `W_DATA_BITWIDTH'b11111_11011110010,
        `W_DATA_BITWIDTH'b11111_11011101011,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b00000_00100001011,
        `W_DATA_BITWIDTH'b00000_00011110000,
        `W_DATA_BITWIDTH'b11111_11011000011,
        `W_DATA_BITWIDTH'b00000_00011010101,
        `W_DATA_BITWIDTH'b00000_00100011101,
        `W_DATA_BITWIDTH'b00000_00011101001,
        `W_DATA_BITWIDTH'b11111_11101111000,
        `W_DATA_BITWIDTH'b00000_00101010111,
        `W_DATA_BITWIDTH'b00000_00010010001,
        `W_DATA_BITWIDTH'b11111_11101011110,
        `W_DATA_BITWIDTH'b00000_00110110001,
        `W_DATA_BITWIDTH'b00000_00100011111,
        `W_DATA_BITWIDTH'b00000_00010001100,
        `W_DATA_BITWIDTH'b00000_01000001001,
        `W_DATA_BITWIDTH'b00000_00010011010,
        `W_DATA_BITWIDTH'b00000_00100011010,
        `W_DATA_BITWIDTH'b00000_00110010110,
        `W_DATA_BITWIDTH'b00000_00010011110,
        `W_DATA_BITWIDTH'b00000_00110111000,
        `W_DATA_BITWIDTH'b00000_00011111101,
        `W_DATA_BITWIDTH'b11111_11001011110,
        `W_DATA_BITWIDTH'b00000_00011111011,
        `W_DATA_BITWIDTH'b11111_11100010100,
        `W_DATA_BITWIDTH'b00000_00011101101,
        `W_DATA_BITWIDTH'b00000_00011010101,
        `W_DATA_BITWIDTH'b00000_00011010101,
        `W_DATA_BITWIDTH'b11111_11100111001,
        `W_DATA_BITWIDTH'b00000_00010100000,
        `W_DATA_BITWIDTH'b11111_11010011010,
        `W_DATA_BITWIDTH'b11111_10111110110,
        `W_DATA_BITWIDTH'b00000_00101110100,
        `W_DATA_BITWIDTH'b00000_00110001101,
        `W_DATA_BITWIDTH'b11111_11001110000,
        `W_DATA_BITWIDTH'b11111_11100101111,
        `W_DATA_BITWIDTH'b11111_11101011011,
        `W_DATA_BITWIDTH'b00000_00010001110,
        `W_DATA_BITWIDTH'b00000_00101110011,
        `W_DATA_BITWIDTH'b11111_11101100111,
        `W_DATA_BITWIDTH'b11111_10101111011,
        `W_DATA_BITWIDTH'b00000_01001101010,
        `W_DATA_BITWIDTH'b00000_00100110000,
        `W_DATA_BITWIDTH'b11111_10001100010,
        `W_DATA_BITWIDTH'b00000_01001110100,
        `W_DATA_BITWIDTH'b00000_00111000100,
        `W_DATA_BITWIDTH'b11111_11011110111,
        `W_DATA_BITWIDTH'b11111_10110100111,
        `W_DATA_BITWIDTH'b00000_00011101011,
        `W_DATA_BITWIDTH'b11111_11000001000,
        `W_DATA_BITWIDTH'b11111_11101001000,
        `W_DATA_BITWIDTH'b00000_00110011101,
        `W_DATA_BITWIDTH'b11111_11010011010,
        `W_DATA_BITWIDTH'b11111_10100100100,
        `W_DATA_BITWIDTH'b00000_00101000100,
        `W_DATA_BITWIDTH'b00000_00110101011,
        `W_DATA_BITWIDTH'b11111_11010111010,
        `W_DATA_BITWIDTH'b11111_11101101000,
        `W_DATA_BITWIDTH'b11111_11101011100,
        `W_DATA_BITWIDTH'b00000_00100010111,
        `W_DATA_BITWIDTH'b00000_00101100010,
        `W_DATA_BITWIDTH'b11111_11000011100,
        `W_DATA_BITWIDTH'b00000_00011001011,
        `W_DATA_BITWIDTH'b11111_11100000011,
        `W_DATA_BITWIDTH'b11111_11011010111,
        `W_DATA_BITWIDTH'b00000_00101111110,
        `W_DATA_BITWIDTH'b00000_00011101001,
        `W_DATA_BITWIDTH'b11111_10011111000,
        `W_DATA_BITWIDTH'b11111_11001001011,
        `W_DATA_BITWIDTH'b00000_00010100101,
        `W_DATA_BITWIDTH'b11111_11011100011,
        `W_DATA_BITWIDTH'b11111_11001001100,
        `W_DATA_BITWIDTH'b11111_11100011000,
        `W_DATA_BITWIDTH'b11111_11001110010,
        `W_DATA_BITWIDTH'b11111_11101110100,
        `W_DATA_BITWIDTH'b00000_00101101000,
        `W_DATA_BITWIDTH'b11111_11001101100,
        `W_DATA_BITWIDTH'b11111_11010110000,
        `W_DATA_BITWIDTH'b11111_11101111001,
        `W_DATA_BITWIDTH'b00000_00011111011,
        `W_DATA_BITWIDTH'b11111_11010010100,
        `W_DATA_BITWIDTH'b00000_00101010000,
        `W_DATA_BITWIDTH'b11111_11100001010,
        `W_DATA_BITWIDTH'b11111_11011110001,
        `W_DATA_BITWIDTH'b00000_00011101010,
        `W_DATA_BITWIDTH'b11111_11101011011,
        `W_DATA_BITWIDTH'b11111_11100101101,
        `W_DATA_BITWIDTH'b11111_11000101000,
        `W_DATA_BITWIDTH'b11111_11100111100,
        `W_DATA_BITWIDTH'b00000_00101001000,
        `W_DATA_BITWIDTH'b00000_00110000010,
        `W_DATA_BITWIDTH'b11111_11010110001,
        `W_DATA_BITWIDTH'b00000_00010110101,
        `W_DATA_BITWIDTH'b11111_11001011100,
        `W_DATA_BITWIDTH'b00000_00011001110,
        `W_DATA_BITWIDTH'b11111_11100010101,
        `W_DATA_BITWIDTH'b11111_11101001101,
        `W_DATA_BITWIDTH'b11111_11011011111,
        `W_DATA_BITWIDTH'b00000_00011110111,
        `W_DATA_BITWIDTH'b11111_11010101110,
        `W_DATA_BITWIDTH'b00000_00010110000,
        `W_DATA_BITWIDTH'b11111_11100100010,
        `W_DATA_BITWIDTH'b00000_00011100100,
        `W_DATA_BITWIDTH'b00000_00100001000,
        `W_DATA_BITWIDTH'b11111_11100100000,
        `W_DATA_BITWIDTH'b00000_00011011100,
        `W_DATA_BITWIDTH'b00000_00101000101,
        `W_DATA_BITWIDTH'b00000_00011000001,
        `W_DATA_BITWIDTH'b00000_00010101110,
        `W_DATA_BITWIDTH'b11111_11100101101,
        `W_DATA_BITWIDTH'b11111_11011111111,
        `W_DATA_BITWIDTH'b00000_00011101001,
        `W_DATA_BITWIDTH'b00000_00010111100,
        `W_DATA_BITWIDTH'b00000_00010101011,
        `W_DATA_BITWIDTH'b00000_00011011100,
        `W_DATA_BITWIDTH'b00000_00010000110,
        `W_DATA_BITWIDTH'b00000_00010010111,
        `W_DATA_BITWIDTH'b00000_00100101011,
        `W_DATA_BITWIDTH'b00000_00101101101,
        `W_DATA_BITWIDTH'b11111_11101110110,
        `W_DATA_BITWIDTH'b11111_10101001100,
        `W_DATA_BITWIDTH'b11111_11100100011,
        `W_DATA_BITWIDTH'b11111_11101000101,
        `W_DATA_BITWIDTH'b00000_00010100011,
        `W_DATA_BITWIDTH'b11111_11101010111,
        `W_DATA_BITWIDTH'b11111_11011111101,
        `W_DATA_BITWIDTH'b11111_11011111010,
        `W_DATA_BITWIDTH'b00000_00100101111,
        `W_DATA_BITWIDTH'b00000_00010000011,
        `W_DATA_BITWIDTH'b00000_00011101111,
        `W_DATA_BITWIDTH'b00000_00010001100,
        `W_DATA_BITWIDTH'b00000_00010001110,
        `W_DATA_BITWIDTH'b11111_11101100001,
        `W_DATA_BITWIDTH'b00000_00010000110,
        `W_DATA_BITWIDTH'b11111_11100110110,
        `W_DATA_BITWIDTH'b00000_00010111011,
        `W_DATA_BITWIDTH'b00000_00010110000,
        `W_DATA_BITWIDTH'b00000_00100000111,
        `W_DATA_BITWIDTH'b00000_00100001111,
        `W_DATA_BITWIDTH'b11111_11011000001,
        `W_DATA_BITWIDTH'b11111_11001100000,
        `W_DATA_BITWIDTH'b11111_11100110110,
        `W_DATA_BITWIDTH'b11111_10110000111,
        `W_DATA_BITWIDTH'b11111_11100101001,
        `W_DATA_BITWIDTH'b11111_11010011101,
        `W_DATA_BITWIDTH'b00000_00101000110,
        `W_DATA_BITWIDTH'b00000_00101100011,
        `W_DATA_BITWIDTH'b00000_00010100101,
        `W_DATA_BITWIDTH'b00000_00101011011,
        `W_DATA_BITWIDTH'b11111_11100011111,
        `W_DATA_BITWIDTH'b11111_11001100010,
        `W_DATA_BITWIDTH'b00000_00100011000,
        `W_DATA_BITWIDTH'b00000_00100010011,
        `W_DATA_BITWIDTH'b11111_11101110011,
        `W_DATA_BITWIDTH'b00000_00011001100,
        `W_DATA_BITWIDTH'b00000_00100111011,
        `W_DATA_BITWIDTH'b11111_11010001011,
        `W_DATA_BITWIDTH'b11111_11100000111,
        `W_DATA_BITWIDTH'b00000_01001000101,
        `W_DATA_BITWIDTH'b11111_11101001111,
        `W_DATA_BITWIDTH'b11111_11010010110,
        `W_DATA_BITWIDTH'b00000_01000111001,
        `W_DATA_BITWIDTH'b00000_00111110000,
        `W_DATA_BITWIDTH'b11111_11101101001,
        `W_DATA_BITWIDTH'b11111_11001101010,
        `W_DATA_BITWIDTH'b11111_11011001000,
        `W_DATA_BITWIDTH'b00000_00011011011,
        `W_DATA_BITWIDTH'b11111_10110110101,
        `W_DATA_BITWIDTH'b11111_11100000000,
        `W_DATA_BITWIDTH'b00000_00010101000,
        `W_DATA_BITWIDTH'b00000_00100000110,
        `W_DATA_BITWIDTH'b00000_01000000111,
        `W_DATA_BITWIDTH'b00000_00100111100,
        `W_DATA_BITWIDTH'b00000_00100111100
    };





// output logic
// logic o_finished_n,


// w_data
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l1_s0_n [0:`W_C_LENGTH_L1_S0-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l1_s1_n [0:`W_C_LENGTH_L1_S1-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l1_s2_n [0:`W_C_LENGTH_L1_S2-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l2_s0_n [0:`W_C_LENGTH_L2_S0-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l2_s1_n [0:`W_C_LENGTH_L2_S1-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l2_s2_n [0:`W_C_LENGTH_L2_S2-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l3_s0_n [0:`W_C_LENGTH_L3_S0-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l3_s1_n [0:`W_C_LENGTH_L3_S1-1];
    logic signed [`W_DATA_BITWIDTH-1 :0] o_w_data_l3_s2_n [0:`W_C_LENGTH_L3_S2-1];

// w_c_idx
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l1_s0_n [0:`W_C_LENGTH_L1_S0-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l1_s1_n [0:`W_C_LENGTH_L1_S1-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l1_s2_n [0:`W_C_LENGTH_L1_S2-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l2_s0_n [0:`W_C_LENGTH_L2_S0-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l2_s1_n [0:`W_C_LENGTH_L2_S1-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l2_s2_n [0:`W_C_LENGTH_L2_S2-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l3_s0_n [0:`W_C_LENGTH_L3_S0-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l3_s1_n [0:`W_C_LENGTH_L3_S1-1];
    logic [`W_C_BITWIDTH-1 :0] o_w_c_idx_l3_s2_n [0:`W_C_LENGTH_L3_S2-1];

// w_r_idx
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l1_s0_n [0:`W_R_LENGTH_L1_S0-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l1_s1_n [0:`W_R_LENGTH_L1_S1-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l1_s2_n [0:`W_R_LENGTH_L1_S2-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l2_s0_n [0:`W_R_LENGTH_L2_S0-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l2_s1_n [0:`W_R_LENGTH_L2_S1-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l2_s2_n [0:`W_R_LENGTH_L2_S2-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l3_s0_n [0:`W_R_LENGTH_L3_S0-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l3_s1_n [0:`W_R_LENGTH_L3_S1-1];
    logic [`W_R_BITWIDTH-1 :0] o_w_r_idx_l3_s2_n [0:`W_R_LENGTH_L3_S2-1];

//  w_k-idx
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l1_s0_n [0:`W_R_LENGTH_L1_S0-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l1_s1_n [0:`W_R_LENGTH_L1_S1-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l1_s2_n [0:`W_R_LENGTH_L1_S2-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l2_s0_n [0:`W_R_LENGTH_L2_S0-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l2_s1_n [0:`W_R_LENGTH_L2_S1-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l2_s2_n [0:`W_R_LENGTH_L2_S2-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l3_s0_n [0:`W_R_LENGTH_L3_S0-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l3_s1_n [0:`W_R_LENGTH_L3_S1-1];
    logic [`W_K_BITWIDTH-1 :0] o_w_k_idx_l3_s2_n [0:`W_R_LENGTH_L3_S2-1];

// w_pos_ptr
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l1_s0_n [0:`W_R_LENGTH_L1_S0-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l1_s1_n [0:`W_R_LENGTH_L1_S1-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l1_s2_n [0:`W_R_LENGTH_L1_S2-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l2_s0_n [0:`W_R_LENGTH_L2_S0-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l2_s1_n [0:`W_R_LENGTH_L2_S1-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l2_s2_n [0:`W_R_LENGTH_L2_S2-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l3_s0_n [0:`W_R_LENGTH_L3_S0-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l3_s1_n [0:`W_R_LENGTH_L3_S1-1];
    logic [`W_POS_PTR_BITWIDTH-1 :0] o_w_pos_ptr_l3_s2_n [0:`W_R_LENGTH_L3_S2-1];



// localparam logic signed [23:0]W_data_l1_s0[6:0] = 
// '{
//     24'b1000_0000_0_1001_000_0010_1100,
//     24'b1001_1000_0_0001_000_0010_1100,
//     24'b0100_0010_0_1110_000_0010_1100,
//     24'b0000_0000_0_0110_000_0010_1100,
//     24'b0000_0000_0_1010_000_0010_1100,
//     24'b1010_1000_0_0010_000_0010_1100,
//     24'b0000_0000_0_1111_000_0010_1100
// };





// =====  logic buffers =====
// assign o_finished = o_finished_r;

// ===== Testing Combinational Blocks =====
always_comb begin 

    // w_data
    for(int k=0; k<`W_C_LENGTH_L1_S0; k=k+1) o_w_data_l1_s0_n[k] = o_w_data_l1_s0[k];
    for(int k=0; k<`W_C_LENGTH_L1_S1; k=k+1) o_w_data_l1_s1_n[k] = o_w_data_l1_s1[k];
    for(int k=0; k<`W_C_LENGTH_L1_S2; k=k+1) o_w_data_l1_s2_n[k] = o_w_data_l1_s2[k];
    for(int k=0; k<`W_C_LENGTH_L2_S0; k=k+1) o_w_data_l2_s0_n[k] = o_w_data_l2_s0[k];
    for(int k=0; k<`W_C_LENGTH_L2_S1; k=k+1) o_w_data_l2_s1_n[k] = o_w_data_l2_s1[k];
    for(int k=0; k<`W_C_LENGTH_L2_S2; k=k+1) o_w_data_l2_s2_n[k] = o_w_data_l2_s2[k];
    for(int k=0; k<`W_C_LENGTH_L3_S0; k=k+1) o_w_data_l3_s0_n[k] = o_w_data_l3_s0[k];
    for(int k=0; k<`W_C_LENGTH_L3_S1; k=k+1) o_w_data_l3_s1_n[k] = o_w_data_l3_s1[k];
    for(int k=0; k<`W_C_LENGTH_L3_S2; k=k+1) o_w_data_l3_s2_n[k] = o_w_data_l3_s2[k];

    // w_c_idx
    for(int k=0; k<`W_C_LENGTH_L1_S0; k=k+1) o_w_c_idx_l1_s0_n[k] = o_w_c_idx_l1_s0[k];
    for(int k=0; k<`W_C_LENGTH_L1_S1; k=k+1) o_w_c_idx_l1_s1_n[k] = o_w_c_idx_l1_s1[k];
    for(int k=0; k<`W_C_LENGTH_L1_S2; k=k+1) o_w_c_idx_l1_s2_n[k] = o_w_c_idx_l1_s2[k];
    for(int k=0; k<`W_C_LENGTH_L2_S0; k=k+1) o_w_c_idx_l2_s0_n[k] = o_w_c_idx_l2_s0[k];
    for(int k=0; k<`W_C_LENGTH_L2_S1; k=k+1) o_w_c_idx_l2_s1_n[k] = o_w_c_idx_l2_s1[k];
    for(int k=0; k<`W_C_LENGTH_L2_S2; k=k+1) o_w_c_idx_l2_s2_n[k] = o_w_c_idx_l2_s2[k];
    for(int k=0; k<`W_C_LENGTH_L3_S0; k=k+1) o_w_c_idx_l3_s0_n[k] = o_w_c_idx_l3_s0[k];
    for(int k=0; k<`W_C_LENGTH_L3_S1; k=k+1) o_w_c_idx_l3_s1_n[k] = o_w_c_idx_l3_s1[k];
    for(int k=0; k<`W_C_LENGTH_L3_S2; k=k+1) o_w_c_idx_l3_s2_n[k] = o_w_c_idx_l3_s2[k];

    // w_r_idx
    for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_r_idx_l1_s0_n[k] = o_w_r_idx_l1_s0[k];
    for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_r_idx_l1_s1_n[k] = o_w_r_idx_l1_s1[k];
    for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_r_idx_l1_s2_n[k] = o_w_r_idx_l1_s2[k];
    for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_r_idx_l2_s0_n[k] = o_w_r_idx_l2_s0[k];
    for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_r_idx_l2_s1_n[k] = o_w_r_idx_l2_s1[k];
    for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_r_idx_l2_s2_n[k] = o_w_r_idx_l2_s2[k];
    for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_r_idx_l3_s0_n[k] = o_w_r_idx_l3_s0[k];
    for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_r_idx_l3_s1_n[k] = o_w_r_idx_l3_s1[k];
    for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_r_idx_l3_s2_n[k] = o_w_r_idx_l3_s2[k];

    // w_k_idx
    for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_k_idx_l1_s0_n[k] = o_w_k_idx_l1_s0[k];
    for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_k_idx_l1_s1_n[k] = o_w_k_idx_l1_s1[k];
    for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_k_idx_l1_s2_n[k] = o_w_k_idx_l1_s2[k];
    for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_k_idx_l2_s0_n[k] = o_w_k_idx_l2_s0[k];
    for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_k_idx_l2_s1_n[k] = o_w_k_idx_l2_s1[k];
    for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_k_idx_l2_s2_n[k] = o_w_k_idx_l2_s2[k];
    for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_k_idx_l3_s0_n[k] = o_w_k_idx_l3_s0[k];
    for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_k_idx_l3_s1_n[k] = o_w_k_idx_l3_s1[k];
    for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_k_idx_l3_s2_n[k] = o_w_k_idx_l3_s2[k];

    // w_posptr
    for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_pos_ptr_l1_s0_n[k] = o_w_pos_ptr_l1_s0[k];
    for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_pos_ptr_l1_s1_n[k] = o_w_pos_ptr_l1_s1[k];
    for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_pos_ptr_l1_s2_n[k] = o_w_pos_ptr_l1_s2[k];
    for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_pos_ptr_l2_s0_n[k] = o_w_pos_ptr_l2_s0[k];
    for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_pos_ptr_l2_s1_n[k] = o_w_pos_ptr_l2_s1[k];
    for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_pos_ptr_l2_s2_n[k] = o_w_pos_ptr_l2_s2[k];
    for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_pos_ptr_l3_s0_n[k] = o_w_pos_ptr_l3_s0[k];
    for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_pos_ptr_l3_s1_n[k] = o_w_pos_ptr_l3_s1[k];
    for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_pos_ptr_l3_s2_n[k] = o_w_pos_ptr_l3_s2[k];
end




// ===== Sequential blocks =====
always_ff @( posedge i_clk or negedge i_rst_n ) begin 
    if(!i_rst_n) begin

        // w_data
        for(int k=0; k<`W_C_LENGTH_L1_S0; k=k+1) o_w_data_l1_s0[k] <= w_data_l1_s0[k];
        for(int k=0; k<`W_C_LENGTH_L1_S1; k=k+1) o_w_data_l1_s1[k] <= w_data_l1_s1[k];
        for(int k=0; k<`W_C_LENGTH_L1_S2; k=k+1) o_w_data_l1_s2[k] <= w_data_l1_s2[k];
        for(int k=0; k<`W_C_LENGTH_L2_S0; k=k+1) o_w_data_l2_s0[k] <= w_data_l2_s0[k];
        for(int k=0; k<`W_C_LENGTH_L2_S1; k=k+1) o_w_data_l2_s1[k] <= w_data_l2_s1[k];
        for(int k=0; k<`W_C_LENGTH_L2_S2; k=k+1) o_w_data_l2_s2[k] <= w_data_l2_s2[k];
        for(int k=0; k<`W_C_LENGTH_L3_S0; k=k+1) o_w_data_l3_s0[k] <= w_data_l3_s0[k];
        for(int k=0; k<`W_C_LENGTH_L3_S1; k=k+1) o_w_data_l3_s1[k] <= w_data_l3_s1[k];
        for(int k=0; k<`W_C_LENGTH_L3_S2; k=k+1) o_w_data_l3_s2[k] <= w_data_l3_s2[k];

        // w_c_idx
        for(int k=0; k<`W_C_LENGTH_L1_S0; k=k+1) o_w_c_idx_l1_s0[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L1_S1; k=k+1) o_w_c_idx_l1_s1[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L1_S2; k=k+1) o_w_c_idx_l1_s2[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L2_S0; k=k+1) o_w_c_idx_l2_s0[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L2_S1; k=k+1) o_w_c_idx_l2_s1[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L2_S2; k=k+1) o_w_c_idx_l2_s2[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L3_S0; k=k+1) o_w_c_idx_l3_s0[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L3_S1; k=k+1) o_w_c_idx_l3_s1[k] <= 0;
        for(int k=0; k<`W_C_LENGTH_L3_S2; k=k+1) o_w_c_idx_l3_s2[k] <= 0;

        // w_r_idx
        for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_r_idx_l1_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_r_idx_l1_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_r_idx_l1_s2[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_r_idx_l2_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_r_idx_l2_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_r_idx_l2_s2[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_r_idx_l3_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_r_idx_l3_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_r_idx_l3_s2[k] <= 0;

        // w_k_idx
        for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_k_idx_l1_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_k_idx_l1_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_k_idx_l1_s2[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_k_idx_l2_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_k_idx_l2_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_k_idx_l2_s2[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_k_idx_l3_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_k_idx_l3_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_k_idx_l3_s2[k] <= 0;

        // w_posptr
        for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_pos_ptr_l1_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_pos_ptr_l1_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_pos_ptr_l1_s2[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_pos_ptr_l2_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_pos_ptr_l2_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_pos_ptr_l2_s2[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_pos_ptr_l3_s0[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_pos_ptr_l3_s1[k] <= 0;
        for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_pos_ptr_l3_s2[k] <= 0;
    end
    else begin

        // w_data
        for(int k=0; k<`W_C_LENGTH_L1_S0; k=k+1) o_w_data_l1_s0[k] <= o_w_data_l1_s0_n[k];
        for(int k=0; k<`W_C_LENGTH_L1_S1; k=k+1) o_w_data_l1_s1[k] <= o_w_data_l1_s1_n[k];
        for(int k=0; k<`W_C_LENGTH_L1_S2; k=k+1) o_w_data_l1_s2[k] <= o_w_data_l1_s2_n[k];
        for(int k=0; k<`W_C_LENGTH_L2_S0; k=k+1) o_w_data_l2_s0[k] <= o_w_data_l2_s0_n[k];
        for(int k=0; k<`W_C_LENGTH_L2_S1; k=k+1) o_w_data_l2_s1[k] <= o_w_data_l2_s1_n[k];
        for(int k=0; k<`W_C_LENGTH_L2_S2; k=k+1) o_w_data_l2_s2[k] <= o_w_data_l2_s2_n[k];
        for(int k=0; k<`W_C_LENGTH_L3_S0; k=k+1) o_w_data_l3_s0[k] <= o_w_data_l3_s0_n[k];
        for(int k=0; k<`W_C_LENGTH_L3_S1; k=k+1) o_w_data_l3_s1[k] <= o_w_data_l3_s1_n[k];
        for(int k=0; k<`W_C_LENGTH_L3_S2; k=k+1) o_w_data_l3_s2[k] <= o_w_data_l3_s2_n[k];

        // w_c_idx
        for(int k=0; k<`W_C_LENGTH_L1_S0; k=k+1) o_w_c_idx_l1_s0[k] <= o_w_c_idx_l1_s0_n[k];
        for(int k=0; k<`W_C_LENGTH_L1_S1; k=k+1) o_w_c_idx_l1_s1[k] <= o_w_c_idx_l1_s1_n[k];
        for(int k=0; k<`W_C_LENGTH_L1_S2; k=k+1) o_w_c_idx_l1_s2[k] <= o_w_c_idx_l1_s2_n[k];
        for(int k=0; k<`W_C_LENGTH_L2_S0; k=k+1) o_w_c_idx_l2_s0[k] <= o_w_c_idx_l2_s0_n[k];
        for(int k=0; k<`W_C_LENGTH_L2_S1; k=k+1) o_w_c_idx_l2_s1[k] <= o_w_c_idx_l2_s1_n[k];
        for(int k=0; k<`W_C_LENGTH_L2_S2; k=k+1) o_w_c_idx_l2_s2[k] <= o_w_c_idx_l2_s2_n[k];
        for(int k=0; k<`W_C_LENGTH_L3_S0; k=k+1) o_w_c_idx_l3_s0[k] <= o_w_c_idx_l3_s0_n[k];
        for(int k=0; k<`W_C_LENGTH_L3_S1; k=k+1) o_w_c_idx_l3_s1[k] <= o_w_c_idx_l3_s1_n[k];
        for(int k=0; k<`W_C_LENGTH_L3_S2; k=k+1) o_w_c_idx_l3_s2[k] <= o_w_c_idx_l3_s2_n[k];

        // w_r_idx
        for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_r_idx_l1_s0[k] <= o_w_r_idx_l1_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_r_idx_l1_s1[k] <= o_w_r_idx_l1_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_r_idx_l1_s2[k] <= o_w_r_idx_l1_s2_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_r_idx_l2_s0[k] <= o_w_r_idx_l2_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_r_idx_l2_s1[k] <= o_w_r_idx_l2_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_r_idx_l2_s2[k] <= o_w_r_idx_l2_s2_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_r_idx_l3_s0[k] <= o_w_r_idx_l3_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_r_idx_l3_s1[k] <= o_w_r_idx_l3_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_r_idx_l3_s2[k] <= o_w_r_idx_l3_s2_n[k];

        // w_k_idx
        for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_k_idx_l1_s0[k] <= o_w_k_idx_l1_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_k_idx_l1_s1[k] <= o_w_k_idx_l1_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_k_idx_l1_s2[k] <= o_w_k_idx_l1_s2_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_k_idx_l2_s0[k] <= o_w_k_idx_l2_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_k_idx_l2_s1[k] <= o_w_k_idx_l2_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_k_idx_l2_s2[k] <= o_w_k_idx_l2_s2_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_k_idx_l3_s0[k] <= o_w_k_idx_l3_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_k_idx_l3_s1[k] <= o_w_k_idx_l3_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_k_idx_l3_s2[k] <= o_w_k_idx_l3_s2_n[k];

        // w_posptr
        for(int k=0; k<`W_R_LENGTH_L1_S0; k=k+1) o_w_pos_ptr_l1_s0[k] <= o_w_pos_ptr_l1_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L1_S1; k=k+1) o_w_pos_ptr_l1_s1[k] <= o_w_pos_ptr_l1_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L1_S2; k=k+1) o_w_pos_ptr_l1_s2[k] <= o_w_pos_ptr_l1_s2_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S0; k=k+1) o_w_pos_ptr_l2_s0[k] <= o_w_pos_ptr_l2_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S1; k=k+1) o_w_pos_ptr_l2_s1[k] <= o_w_pos_ptr_l2_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L2_S2; k=k+1) o_w_pos_ptr_l2_s2[k] <= o_w_pos_ptr_l2_s2_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S0; k=k+1) o_w_pos_ptr_l3_s0[k] <= o_w_pos_ptr_l3_s0_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S1; k=k+1) o_w_pos_ptr_l3_s1[k] <= o_w_pos_ptr_l3_s1_n[k];
        for(int k=0; k<`W_R_LENGTH_L3_S2; k=k+1) o_w_pos_ptr_l3_s2[k] <= o_w_pos_ptr_l3_s2_n[k];
    end
end
endmodule
