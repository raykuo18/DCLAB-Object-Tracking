`timescale 1us/1us


// --------------------- `define for WMem ------------------------
    `define W_DATA_BITWIDTH    16
    `define W_C_BITWIDTH       5   // log2(# Channel)
    `define W_R_BITWIDTH       2 
    `define W_K_BITWIDTH       5 
    `define W_POS_PTR_BITWIDTH 11 

    `define W_C_LENGTH_L1_S0  123
    `define W_R_LENGTH_L1_S0  48
    `define W_C_LENGTH_L1_S1  130
    `define W_R_LENGTH_L1_S1  48
    `define W_C_LENGTH_L1_S2  124
    `define W_R_LENGTH_L1_S2  48

    `define W_C_LENGTH_L2_S0  474
    `define W_R_LENGTH_L2_S0  48
    `define W_C_LENGTH_L2_S1  460
    `define W_R_LENGTH_L2_S1  48
    `define W_C_LENGTH_L2_S2  446
    `define W_R_LENGTH_L2_S2  48

    `define W_C_LENGTH        474 // max of C_LENGTH
    `define W_R_LENGTH        48  // max of R_LENGTH


// --------------------- `define for IA ------------------------
    `define IA_DATA_BITWIDTH    16
    `define IA_C_BITWIDTH       5   // log2(# Channel)
    `define IA_CHANNEL 8
    `define IA_ROW 16
    `define IA_COL 16





module tb_PE_TEMP;
	localparam CLK = 10;
	localparam HCLK = CLK/2;

	logic rst, clk;
	initial clk = 0;
	always #HCLK clk = ~clk;



      // ========================== Parameters definition ==================================

        // ----- WMem --------
            // w_data
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
                '{
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b1111110111110001,
                    `W_DATA_BITWIDTH'b0000000010111001,
                    `W_DATA_BITWIDTH'b1111111001001000,
                    `W_DATA_BITWIDTH'b1111111100101100,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000001011101001,
                    `W_DATA_BITWIDTH'b0000001110000101,
                    `W_DATA_BITWIDTH'b1111100101001100,
                    `W_DATA_BITWIDTH'b1111101000011010,
                    `W_DATA_BITWIDTH'b0000001000111111,
                    `W_DATA_BITWIDTH'b1111011110101000,
                    `W_DATA_BITWIDTH'b1111111011101100,
                    `W_DATA_BITWIDTH'b0000110100100001,
                    `W_DATA_BITWIDTH'b0000011110000000,
                    `W_DATA_BITWIDTH'b1111011101111100,
                    `W_DATA_BITWIDTH'b0000101111111011,
                    `W_DATA_BITWIDTH'b1111110110101010,
                    `W_DATA_BITWIDTH'b0000010000001010,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b1111001101110010,
                    `W_DATA_BITWIDTH'b0000101101101000,
                    `W_DATA_BITWIDTH'b0000001101100100,
                    `W_DATA_BITWIDTH'b0000100001011110,
                    `W_DATA_BITWIDTH'b1111101101101010,
                    `W_DATA_BITWIDTH'b0000010110010101,
                    `W_DATA_BITWIDTH'b0000100011000111,
                    `W_DATA_BITWIDTH'b1111111001000000,
                    `W_DATA_BITWIDTH'b1111101000010001,
                    `W_DATA_BITWIDTH'b0000000111110100,
                    `W_DATA_BITWIDTH'b0000001111001101,
                    `W_DATA_BITWIDTH'b0000100001011110,
                    `W_DATA_BITWIDTH'b0000010110100100,
                    `W_DATA_BITWIDTH'b0000001001101110,
                    `W_DATA_BITWIDTH'b1111110000000001,
                    `W_DATA_BITWIDTH'b1111100111111011,
                    `W_DATA_BITWIDTH'b1111101010101100,
                    `W_DATA_BITWIDTH'b1111011110100100,
                    `W_DATA_BITWIDTH'b0000011011011001,
                    `W_DATA_BITWIDTH'b1111101111111110,
                    `W_DATA_BITWIDTH'b0000010000110000,
                    `W_DATA_BITWIDTH'b1111110110111010,
                    `W_DATA_BITWIDTH'b1111100011101101,
                    `W_DATA_BITWIDTH'b1111110010001101,
                    `W_DATA_BITWIDTH'b0000001110100011,
                    `W_DATA_BITWIDTH'b0000011111010101,
                    `W_DATA_BITWIDTH'b1111101110111101,
                    `W_DATA_BITWIDTH'b0000010101111100,
                    `W_DATA_BITWIDTH'b0000001011110110,
                    `W_DATA_BITWIDTH'b0000010010100011,
                    `W_DATA_BITWIDTH'b0000000100100010,
                    `W_DATA_BITWIDTH'b0000010110111000,
                    `W_DATA_BITWIDTH'b0000000100101001,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000111000001,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111001101111,
                    `W_DATA_BITWIDTH'b1111111000010110,
                    `W_DATA_BITWIDTH'b0000000111101010,
                    `W_DATA_BITWIDTH'b0000000111001111,
                    `W_DATA_BITWIDTH'b1111110101100100,
                    `W_DATA_BITWIDTH'b0000010001001100,
                    `W_DATA_BITWIDTH'b0000010010000011,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000100101011,
                    `W_DATA_BITWIDTH'b0000001001100011,
                    `W_DATA_BITWIDTH'b1111101111010111,
                    `W_DATA_BITWIDTH'b1111101010110111,
                    `W_DATA_BITWIDTH'b0000001111100111,
                    `W_DATA_BITWIDTH'b0000001101000010,
                    `W_DATA_BITWIDTH'b1111101110111001,
                    `W_DATA_BITWIDTH'b0000010010101110,
                    `W_DATA_BITWIDTH'b0000001111100110,
                    `W_DATA_BITWIDTH'b0000010010010110,
                    `W_DATA_BITWIDTH'b1111110100101101,
                    `W_DATA_BITWIDTH'b1111111011010101,
                    `W_DATA_BITWIDTH'b1111110100001000,
                    `W_DATA_BITWIDTH'b1111111011001011,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111010100111,
                    `W_DATA_BITWIDTH'b1111111001011111,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111110101010000,
                    `W_DATA_BITWIDTH'b1111111001001110,
                    `W_DATA_BITWIDTH'b1111101010011110,
                    `W_DATA_BITWIDTH'b1111100100101111,
                    `W_DATA_BITWIDTH'b1111110010101000,
                    `W_DATA_BITWIDTH'b1111010110111011,
                    `W_DATA_BITWIDTH'b0000001011110000,
                    `W_DATA_BITWIDTH'b1111110010011011,
                    `W_DATA_BITWIDTH'b0000000111101001,
                    `W_DATA_BITWIDTH'b0000001101010010,
                    `W_DATA_BITWIDTH'b0000000010011101,
                    `W_DATA_BITWIDTH'b1111111000010111,
                    `W_DATA_BITWIDTH'b0000011110111111,
                    `W_DATA_BITWIDTH'b0000100010111000,
                    `W_DATA_BITWIDTH'b0000001000011010,
                    `W_DATA_BITWIDTH'b1111100110001010,
                    `W_DATA_BITWIDTH'b1111110011110100,
                    `W_DATA_BITWIDTH'b1111101011111011,
                    `W_DATA_BITWIDTH'b0000001011001011,
                    `W_DATA_BITWIDTH'b0000001000110010,
                    `W_DATA_BITWIDTH'b1111110010001011,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b1111111101111110,
                    `W_DATA_BITWIDTH'b0000001001111101,
                    `W_DATA_BITWIDTH'b0000001000001111,
                    `W_DATA_BITWIDTH'b1111110111000001,
                    `W_DATA_BITWIDTH'b1111101000000010,
                    `W_DATA_BITWIDTH'b0000010000001111,
                    `W_DATA_BITWIDTH'b1111110101010001,
                    `W_DATA_BITWIDTH'b0000000101110110,
                    `W_DATA_BITWIDTH'b0000001100010100,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b0000000110000101,
                    `W_DATA_BITWIDTH'b1111111100111100,
                    `W_DATA_BITWIDTH'b0000001000011100,
                    `W_DATA_BITWIDTH'b0000001000110011,
                    `W_DATA_BITWIDTH'b0000000110011001,
                    `W_DATA_BITWIDTH'b0000000101111100,
                    `W_DATA_BITWIDTH'b0000001001100000,
                    `W_DATA_BITWIDTH'b1111110110110110,
                    `W_DATA_BITWIDTH'b1111110110110110
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000101011111,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b0000000111100111,
                    `W_DATA_BITWIDTH'b0000000100101110,
                    `W_DATA_BITWIDTH'b0000001000110010,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b1111110111110110,
                    `W_DATA_BITWIDTH'b1111100111000001,
                    `W_DATA_BITWIDTH'b1111110111010101,
                    `W_DATA_BITWIDTH'b1111110000111010,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b0000000011011000,
                    `W_DATA_BITWIDTH'b1111111010010100,
                    `W_DATA_BITWIDTH'b0000000101001111,
                    `W_DATA_BITWIDTH'b1111101100011101,
                    `W_DATA_BITWIDTH'b0000010110011010,
                    `W_DATA_BITWIDTH'b1111110100111010,
                    `W_DATA_BITWIDTH'b1111100010111110,
                    `W_DATA_BITWIDTH'b1111011101011101,
                    `W_DATA_BITWIDTH'b1111011000001011,
                    `W_DATA_BITWIDTH'b1111110101001011,
                    `W_DATA_BITWIDTH'b0000010111101111,
                    `W_DATA_BITWIDTH'b1111111000000100,
                    `W_DATA_BITWIDTH'b0000101110010000,
                    `W_DATA_BITWIDTH'b1111011100111010,
                    `W_DATA_BITWIDTH'b0000001101111000,
                    `W_DATA_BITWIDTH'b1111101010101101,
                    `W_DATA_BITWIDTH'b0000100000101000,
                    `W_DATA_BITWIDTH'b0000101110110101,
                    `W_DATA_BITWIDTH'b1111101100111000,
                    `W_DATA_BITWIDTH'b1111101100011100,
                    `W_DATA_BITWIDTH'b1111011100100010,
                    `W_DATA_BITWIDTH'b0000100000110000,
                    `W_DATA_BITWIDTH'b0000011110000000,
                    `W_DATA_BITWIDTH'b0000011000010101,
                    `W_DATA_BITWIDTH'b0000001010000011,
                    `W_DATA_BITWIDTH'b0000010000010000,
                    `W_DATA_BITWIDTH'b0000000011111110,
                    `W_DATA_BITWIDTH'b1111101100111110,
                    `W_DATA_BITWIDTH'b1111101110110110,
                    `W_DATA_BITWIDTH'b0000001000100110,
                    `W_DATA_BITWIDTH'b0000010011101111,
                    `W_DATA_BITWIDTH'b0000001010110001,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b1111100011110100,
                    `W_DATA_BITWIDTH'b1111100110101001,
                    `W_DATA_BITWIDTH'b0000011101011110,
                    `W_DATA_BITWIDTH'b1111111011101000,
                    `W_DATA_BITWIDTH'b0000001110110001,
                    `W_DATA_BITWIDTH'b0000001101001111,
                    `W_DATA_BITWIDTH'b0000001110100111,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b1111101000011110,
                    `W_DATA_BITWIDTH'b1111100110000110,
                    `W_DATA_BITWIDTH'b0000000111110100,
                    `W_DATA_BITWIDTH'b1111101011101001,
                    `W_DATA_BITWIDTH'b1111111011010000,
                    `W_DATA_BITWIDTH'b0000011100111011,
                    `W_DATA_BITWIDTH'b1111111001010001,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000100001001,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b1111111010010000,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000110101011,
                    `W_DATA_BITWIDTH'b0000000011001110,
                    `W_DATA_BITWIDTH'b0000001011100010,
                    `W_DATA_BITWIDTH'b1111111001100000,
                    `W_DATA_BITWIDTH'b0000010000010010,
                    `W_DATA_BITWIDTH'b0000000100000100,
                    `W_DATA_BITWIDTH'b1111111011101001,
                    `W_DATA_BITWIDTH'b1111101101101001,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111111100100110,
                    `W_DATA_BITWIDTH'b1111110011011001,
                    `W_DATA_BITWIDTH'b1111110011110101,
                    `W_DATA_BITWIDTH'b0000000110111011,
                    `W_DATA_BITWIDTH'b0000001000110011,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b0000010010110111,
                    `W_DATA_BITWIDTH'b0000001000010010,
                    `W_DATA_BITWIDTH'b0000001111100010,
                    `W_DATA_BITWIDTH'b1111101110000101,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b0000000100011110,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b1111101111111100,
                    `W_DATA_BITWIDTH'b0000100011111111,
                    `W_DATA_BITWIDTH'b0000001001011111,
                    `W_DATA_BITWIDTH'b1111011100110011,
                    `W_DATA_BITWIDTH'b0000000101111010,
                    `W_DATA_BITWIDTH'b0000100001010011,
                    `W_DATA_BITWIDTH'b0000100100011011,
                    `W_DATA_BITWIDTH'b1111100011111100,
                    `W_DATA_BITWIDTH'b0000000011100010,
                    `W_DATA_BITWIDTH'b0000000110001010,
                    `W_DATA_BITWIDTH'b0000000101101101,
                    `W_DATA_BITWIDTH'b0000000100110111,
                    `W_DATA_BITWIDTH'b1111110000110011,
                    `W_DATA_BITWIDTH'b1111110011001100,
                    `W_DATA_BITWIDTH'b0000010011110100,
                    `W_DATA_BITWIDTH'b1111100001111001,
                    `W_DATA_BITWIDTH'b1111101011000000,
                    `W_DATA_BITWIDTH'b0000011000110100,
                    `W_DATA_BITWIDTH'b1111111000010010,
                    `W_DATA_BITWIDTH'b1111110101110110,
                    `W_DATA_BITWIDTH'b1111110000001110,
                    `W_DATA_BITWIDTH'b1111110101100100,
                    `W_DATA_BITWIDTH'b0000001110111111,
                    `W_DATA_BITWIDTH'b1111111101110011,
                    `W_DATA_BITWIDTH'b0000000111101110,
                    `W_DATA_BITWIDTH'b0000001100100011,
                    `W_DATA_BITWIDTH'b1111110110110100,
                    `W_DATA_BITWIDTH'b1111111100110101,
                    `W_DATA_BITWIDTH'b0000000111111110,
                    `W_DATA_BITWIDTH'b0000001101111010,
                    `W_DATA_BITWIDTH'b1111111000111010,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b1111110010000001,
                    `W_DATA_BITWIDTH'b1111110000111011,
                    `W_DATA_BITWIDTH'b1111110110111010,
                    `W_DATA_BITWIDTH'b1111111001000010,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b1111110111110111,
                    `W_DATA_BITWIDTH'b0000000111000111,
                    `W_DATA_BITWIDTH'b0000001011100000,
                    `W_DATA_BITWIDTH'b0000000101101011,
                    `W_DATA_BITWIDTH'b0000000101101011
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b1111111001101101,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000101101111,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b0000000110001110,
                    `W_DATA_BITWIDTH'b0000000111000011,
                    `W_DATA_BITWIDTH'b0000000100111000,
                    `W_DATA_BITWIDTH'b0000001010100011,
                    `W_DATA_BITWIDTH'b0000011001010111,
                    `W_DATA_BITWIDTH'b0000010111100000,
                    `W_DATA_BITWIDTH'b1111110101010110,
                    `W_DATA_BITWIDTH'b0000001110110110,
                    `W_DATA_BITWIDTH'b0000010000001100,
                    `W_DATA_BITWIDTH'b0000011101011110,
                    `W_DATA_BITWIDTH'b0000100011000010,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b0000010110101000,
                    `W_DATA_BITWIDTH'b1111110111000001,
                    `W_DATA_BITWIDTH'b1111101101110010,
                    `W_DATA_BITWIDTH'b1111100001100100,
                    `W_DATA_BITWIDTH'b1111011100010000,
                    `W_DATA_BITWIDTH'b0000001010010010,
                    `W_DATA_BITWIDTH'b0000100010011111,
                    `W_DATA_BITWIDTH'b1111111001101100,
                    `W_DATA_BITWIDTH'b1111100000100001,
                    `W_DATA_BITWIDTH'b1111110001100011,
                    `W_DATA_BITWIDTH'b1111110101110110,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b1111011101000001,
                    `W_DATA_BITWIDTH'b1111011110011101,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b0000001110110100,
                    `W_DATA_BITWIDTH'b1111101101011100,
                    `W_DATA_BITWIDTH'b0000000110010011,
                    `W_DATA_BITWIDTH'b1111101000101111,
                    `W_DATA_BITWIDTH'b1111111001100001,
                    `W_DATA_BITWIDTH'b1111110000101001,
                    `W_DATA_BITWIDTH'b1111101101110000,
                    `W_DATA_BITWIDTH'b0000001101010011,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000010011110101,
                    `W_DATA_BITWIDTH'b1111100010100000,
                    `W_DATA_BITWIDTH'b1111011000000110,
                    `W_DATA_BITWIDTH'b1111101001101111,
                    `W_DATA_BITWIDTH'b1111110101000000,
                    `W_DATA_BITWIDTH'b0000001011000000,
                    `W_DATA_BITWIDTH'b0000011010001000,
                    `W_DATA_BITWIDTH'b0000001000110001,
                    `W_DATA_BITWIDTH'b0000010111001000,
                    `W_DATA_BITWIDTH'b1111101010011000,
                    `W_DATA_BITWIDTH'b1111100001101011,
                    `W_DATA_BITWIDTH'b1111111011001100,
                    `W_DATA_BITWIDTH'b1111100010111100,
                    `W_DATA_BITWIDTH'b0000001110101000,
                    `W_DATA_BITWIDTH'b0000000100011011,
                    `W_DATA_BITWIDTH'b0000011111001100,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b0000000101100011,
                    `W_DATA_BITWIDTH'b1111111011001101,
                    `W_DATA_BITWIDTH'b0000001001000110,
                    `W_DATA_BITWIDTH'b0000001001000011,
                    `W_DATA_BITWIDTH'b1111111011101110,
                    `W_DATA_BITWIDTH'b0000001110000101,
                    `W_DATA_BITWIDTH'b0000001110011101,
                    `W_DATA_BITWIDTH'b1111111000001111,
                    `W_DATA_BITWIDTH'b0000001011110001,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b0000000100100001,
                    `W_DATA_BITWIDTH'b0000001011111111,
                    `W_DATA_BITWIDTH'b1111110101010110,
                    `W_DATA_BITWIDTH'b1111111011100001,
                    `W_DATA_BITWIDTH'b1111101101010001,
                    `W_DATA_BITWIDTH'b1111110001110111,
                    `W_DATA_BITWIDTH'b0000001010111101,
                    `W_DATA_BITWIDTH'b1111110001101001,
                    `W_DATA_BITWIDTH'b0000001010100110,
                    `W_DATA_BITWIDTH'b0000001101010001,
                    `W_DATA_BITWIDTH'b1111110001001111,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b1111111011100110,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b0000000101000111,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b0000010111010101,
                    `W_DATA_BITWIDTH'b0000011011111100,
                    `W_DATA_BITWIDTH'b0000011010010110,
                    `W_DATA_BITWIDTH'b0000001000100010,
                    `W_DATA_BITWIDTH'b1111101010000010,
                    `W_DATA_BITWIDTH'b1111111000101001,
                    `W_DATA_BITWIDTH'b1111110110010100,
                    `W_DATA_BITWIDTH'b0000000111011110,
                    `W_DATA_BITWIDTH'b1111101011011110,
                    `W_DATA_BITWIDTH'b0000011111111101,
                    `W_DATA_BITWIDTH'b1111011101110110,
                    `W_DATA_BITWIDTH'b1111110111011101,
                    `W_DATA_BITWIDTH'b1111111000101110,
                    `W_DATA_BITWIDTH'b0000010011001111,
                    `W_DATA_BITWIDTH'b0000001010011000,
                    `W_DATA_BITWIDTH'b1111101011100110,
                    `W_DATA_BITWIDTH'b1111111000011100,
                    `W_DATA_BITWIDTH'b1111111000010110,
                    `W_DATA_BITWIDTH'b1111110101011010,
                    `W_DATA_BITWIDTH'b1111110101001001,
                    `W_DATA_BITWIDTH'b1111111001100010,
                    `W_DATA_BITWIDTH'b0000000110110101,
                    `W_DATA_BITWIDTH'b0000000110111010,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b0000001011100010,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b0000001010000000,
                    `W_DATA_BITWIDTH'b1111111001011011,
                    `W_DATA_BITWIDTH'b1111111011011111,
                    `W_DATA_BITWIDTH'b1111110001101000,
                    `W_DATA_BITWIDTH'b1111110111010101,
                    `W_DATA_BITWIDTH'b1111111010100010,
                    `W_DATA_BITWIDTH'b1111111001011001,
                    `W_DATA_BITWIDTH'b1111111001111110,
                    `W_DATA_BITWIDTH'b0000001010101001,
                    `W_DATA_BITWIDTH'b1111111001011110,
                    `W_DATA_BITWIDTH'b0000000100010001,
                    `W_DATA_BITWIDTH'b1111111000010110,
                    `W_DATA_BITWIDTH'b1111111000010110
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111111101101010,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111001010010,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b0000000010011101,
                    `W_DATA_BITWIDTH'b1111111011010101,
                    `W_DATA_BITWIDTH'b0000000011011001,
                    `W_DATA_BITWIDTH'b0000000100110100,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000010010010,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b0000000110001101,
                    `W_DATA_BITWIDTH'b1111111010111110,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b1111111101001111,
                    `W_DATA_BITWIDTH'b0000000101001001,
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b0000000010001000,
                    `W_DATA_BITWIDTH'b1111111101001110,
                    `W_DATA_BITWIDTH'b1111111100000100,
                    `W_DATA_BITWIDTH'b0000000010111100,
                    `W_DATA_BITWIDTH'b0000000011101000,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b1111111011100111,
                    `W_DATA_BITWIDTH'b1111111101101001,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111100001000,
                    `W_DATA_BITWIDTH'b0000000011000010,
                    `W_DATA_BITWIDTH'b0000000010100100,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b1111111011000111,
                    `W_DATA_BITWIDTH'b0000000011000000,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b1111111001110100,
                    `W_DATA_BITWIDTH'b1111111001000101,
                    `W_DATA_BITWIDTH'b0000000100111001,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b0000000110001111,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b0000000101100010,
                    `W_DATA_BITWIDTH'b1111111100001101,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111011010110,
                    `W_DATA_BITWIDTH'b0000000011011101,
                    `W_DATA_BITWIDTH'b1111110111000000,
                    `W_DATA_BITWIDTH'b1111111001011011,
                    `W_DATA_BITWIDTH'b1111111000101101,
                    `W_DATA_BITWIDTH'b0000000100101110,
                    `W_DATA_BITWIDTH'b0000000011100011,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111110111110011,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b1111111101011101,
                    `W_DATA_BITWIDTH'b0000000100010011,
                    `W_DATA_BITWIDTH'b1111111011011000,
                    `W_DATA_BITWIDTH'b1111111101000011,
                    `W_DATA_BITWIDTH'b1111111101000110,
                    `W_DATA_BITWIDTH'b0000000100010110,
                    `W_DATA_BITWIDTH'b0000000011100001,
                    `W_DATA_BITWIDTH'b1111111011011010,
                    `W_DATA_BITWIDTH'b1111110111011001,
                    `W_DATA_BITWIDTH'b1111111010110110,
                    `W_DATA_BITWIDTH'b1111111011001010,
                    `W_DATA_BITWIDTH'b0000000100001011,
                    `W_DATA_BITWIDTH'b0000000010010100,
                    `W_DATA_BITWIDTH'b1111111011001110,
                    `W_DATA_BITWIDTH'b1111111001100010,
                    `W_DATA_BITWIDTH'b0000000010100101,
                    `W_DATA_BITWIDTH'b1111111010101110,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b1111111010101000,
                    `W_DATA_BITWIDTH'b1111111100111001,
                    `W_DATA_BITWIDTH'b1111111010110010,
                    `W_DATA_BITWIDTH'b0000000010110101,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111100011100,
                    `W_DATA_BITWIDTH'b1111110110001010,
                    `W_DATA_BITWIDTH'b0000000010110111,
                    `W_DATA_BITWIDTH'b0000000111001000,
                    `W_DATA_BITWIDTH'b0000000100101101,
                    `W_DATA_BITWIDTH'b1111111010111001,
                    `W_DATA_BITWIDTH'b0000000011001101,
                    `W_DATA_BITWIDTH'b1111110001110111,
                    `W_DATA_BITWIDTH'b1111111000100001,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b1111110100001001,
                    `W_DATA_BITWIDTH'b1111111010010111,
                    `W_DATA_BITWIDTH'b1111110111001110,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b1111111001001100,
                    `W_DATA_BITWIDTH'b1111110110100001,
                    `W_DATA_BITWIDTH'b1111111011010010,
                    `W_DATA_BITWIDTH'b0000000101110000,
                    `W_DATA_BITWIDTH'b1111111010111010,
                    `W_DATA_BITWIDTH'b1111111011101010,
                    `W_DATA_BITWIDTH'b1111111010100011,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111100100101,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b1111111011011011,
                    `W_DATA_BITWIDTH'b0000000100110100,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b0000000011010111,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b1111111101100000,
                    `W_DATA_BITWIDTH'b0000000010110010,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b0000000100101110,
                    `W_DATA_BITWIDTH'b0000000010100000,
                    `W_DATA_BITWIDTH'b1111111010010101,
                    `W_DATA_BITWIDTH'b1111111101001100,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b1111111010110101,
                    `W_DATA_BITWIDTH'b1111111101111100,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b1111111100110111,
                    `W_DATA_BITWIDTH'b1111111011011100,
                    `W_DATA_BITWIDTH'b1111111100001011,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111100101110,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b1111111011110000,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b0000000100100101,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b1111111010100010,
                    `W_DATA_BITWIDTH'b1111111010110000,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b0000000011010000,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b0000000011000010,
                    `W_DATA_BITWIDTH'b0000000100001101,
                    `W_DATA_BITWIDTH'b0000000011101101,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b1111111011101101,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b1111111101011110,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b0000000101001001,
                    `W_DATA_BITWIDTH'b0000000011000000,
                    `W_DATA_BITWIDTH'b0000000101110110,
                    `W_DATA_BITWIDTH'b0000000010110110,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b0000000011010011,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111111100100010,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000011100001,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b1111111101001001,
                    `W_DATA_BITWIDTH'b1111111101010001,
                    `W_DATA_BITWIDTH'b1111111101100101,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111100001011,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000011100011,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b1111111010101110,
                    `W_DATA_BITWIDTH'b1111111011000011,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b1111111011010011,
                    `W_DATA_BITWIDTH'b1111111101000000,
                    `W_DATA_BITWIDTH'b1111111001111100,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b0000000011101000,
                    `W_DATA_BITWIDTH'b1111111101101111,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b0000000010111001,
                    `W_DATA_BITWIDTH'b1111111101101011,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000100010010,
                    `W_DATA_BITWIDTH'b0000000100110100,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b1111111010110110,
                    `W_DATA_BITWIDTH'b1111111100111110,
                    `W_DATA_BITWIDTH'b0000000100001010,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b0000000101111001,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111011101110,
                    `W_DATA_BITWIDTH'b0000000101111101,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111010100011,
                    `W_DATA_BITWIDTH'b0000000100100011,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b1111110110111010,
                    `W_DATA_BITWIDTH'b1111111101000110,
                    `W_DATA_BITWIDTH'b1111111011001000,
                    `W_DATA_BITWIDTH'b0000000011010001,
                    `W_DATA_BITWIDTH'b1111110001011000,
                    `W_DATA_BITWIDTH'b1111111100000100,
                    `W_DATA_BITWIDTH'b0000000111001101,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b0000000101001011,
                    `W_DATA_BITWIDTH'b0000000110110111,
                    `W_DATA_BITWIDTH'b1111110101001010,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000001000010101,
                    `W_DATA_BITWIDTH'b1111111001010010,
                    `W_DATA_BITWIDTH'b0000000110001000,
                    `W_DATA_BITWIDTH'b0000000011100110,
                    `W_DATA_BITWIDTH'b1111110111000110,
                    `W_DATA_BITWIDTH'b1111111001101001,
                    `W_DATA_BITWIDTH'b1111111001110011,
                    `W_DATA_BITWIDTH'b1111111101001010,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b0000000101010010,
                    `W_DATA_BITWIDTH'b0000000100101000,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b1111111001111100,
                    `W_DATA_BITWIDTH'b1111111100000011,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b0000000110001101,
                    `W_DATA_BITWIDTH'b1111111101001011,
                    `W_DATA_BITWIDTH'b1111111010111110,
                    `W_DATA_BITWIDTH'b1111111001100101,
                    `W_DATA_BITWIDTH'b0000001000110111,
                    `W_DATA_BITWIDTH'b1111111000100010,
                    `W_DATA_BITWIDTH'b1111111100011001,
                    `W_DATA_BITWIDTH'b0000001001000111,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b1111111101111100,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111100101010,
                    `W_DATA_BITWIDTH'b0000000010010100,
                    `W_DATA_BITWIDTH'b1111111100101010,
                    `W_DATA_BITWIDTH'b1111111101010010,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111111101011100,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b1111111100010100,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b1111111011001110,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000100001101,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b1111111101011100,
                    `W_DATA_BITWIDTH'b0000000101100010,
                    `W_DATA_BITWIDTH'b0000000011001001,
                    `W_DATA_BITWIDTH'b1111111011100101,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000011100010,
                    `W_DATA_BITWIDTH'b0000000100011100,
                    `W_DATA_BITWIDTH'b1111111011100111,
                    `W_DATA_BITWIDTH'b0000000110000011,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b1111111011110010,
                    `W_DATA_BITWIDTH'b1111111100101110,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b1111111000010001,
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b1111111011100000,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b1111111100100100,
                    `W_DATA_BITWIDTH'b1111111101101110,
                    `W_DATA_BITWIDTH'b1111111101101100,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111001010001,
                    `W_DATA_BITWIDTH'b1111111101000010,
                    `W_DATA_BITWIDTH'b1111111011111100,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b1111111010111111,
                    `W_DATA_BITWIDTH'b0000000010001010,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b1111111000101010,
                    `W_DATA_BITWIDTH'b0000000100101101,
                    `W_DATA_BITWIDTH'b0000001001100010,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000001010100001,
                    `W_DATA_BITWIDTH'b0000000011001010,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b0000000110001110,
                    `W_DATA_BITWIDTH'b1111111100100001,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b1111111010101101,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000100011010,
                    `W_DATA_BITWIDTH'b1111111100110011,
                    `W_DATA_BITWIDTH'b0000000110101000,
                    `W_DATA_BITWIDTH'b0000000011000000,
                    `W_DATA_BITWIDTH'b0000000111011000,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b0000000111100110,
                    `W_DATA_BITWIDTH'b1111111011111101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000110011101,
                    `W_DATA_BITWIDTH'b1111111101111011,
                    `W_DATA_BITWIDTH'b1111111000111001,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b1111111001001001,
                    `W_DATA_BITWIDTH'b0000000111111000,
                    `W_DATA_BITWIDTH'b1111111001111011,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b1111111011010010,
                    `W_DATA_BITWIDTH'b1111111000011001,
                    `W_DATA_BITWIDTH'b0000000010001010,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111111010000011,
                    `W_DATA_BITWIDTH'b0000000011000110,
                    `W_DATA_BITWIDTH'b1111111001111010,
                    `W_DATA_BITWIDTH'b1111110111011001,
                    `W_DATA_BITWIDTH'b1111111101010001,
                    `W_DATA_BITWIDTH'b1111111001110011,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b0000000101101111,
                    `W_DATA_BITWIDTH'b0000000101011111,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b1111111101110011,
                    `W_DATA_BITWIDTH'b1111111101100010,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111110111100100,
                    `W_DATA_BITWIDTH'b1111111101011111,
                    `W_DATA_BITWIDTH'b0000000011100101,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b1111110110010110,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b0000000110001000,
                    `W_DATA_BITWIDTH'b1111111011101011,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b1111111010001111,
                    `W_DATA_BITWIDTH'b0000000110010101,
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b0000000100000000,
                    `W_DATA_BITWIDTH'b1111111001010000,
                    `W_DATA_BITWIDTH'b0000000011111101,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b0000000010011100,
                    `W_DATA_BITWIDTH'b1111111101111011,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111101001010,
                    `W_DATA_BITWIDTH'b0000000011110101,
                    `W_DATA_BITWIDTH'b0000000100111110,
                    `W_DATA_BITWIDTH'b0000000100011011,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b1111111100110000,
                    `W_DATA_BITWIDTH'b1111111001100110,
                    `W_DATA_BITWIDTH'b0000000011101101,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111001111101,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b1111111010011000,
                    `W_DATA_BITWIDTH'b0000000011001001,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000010011010,
                    `W_DATA_BITWIDTH'b0000000100010001,
                    `W_DATA_BITWIDTH'b1111111011011011,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111011011001,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b1111111011100111,
                    `W_DATA_BITWIDTH'b0000000011111110,
                    `W_DATA_BITWIDTH'b0000000100000100,
                    `W_DATA_BITWIDTH'b0000000010100100,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000011110100,
                    `W_DATA_BITWIDTH'b0000000010010000,
                    `W_DATA_BITWIDTH'b0000000010111000,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b0000000010001010,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b0000000010011100,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b1111110111010111,
                    `W_DATA_BITWIDTH'b1111111001100011,
                    `W_DATA_BITWIDTH'b1111110111111111,
                    `W_DATA_BITWIDTH'b1111110110100011,
                    `W_DATA_BITWIDTH'b0000000010110110,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000101110000,
                    `W_DATA_BITWIDTH'b1111111010110011,
                    `W_DATA_BITWIDTH'b1111111101100010,
                    `W_DATA_BITWIDTH'b1111110111001110,
                    `W_DATA_BITWIDTH'b1111110001110100,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111110110011011,
                    `W_DATA_BITWIDTH'b1111111011111001,
                    `W_DATA_BITWIDTH'b1111111011111000,
                    `W_DATA_BITWIDTH'b0000000100011100,
                    `W_DATA_BITWIDTH'b1111111000001101,
                    `W_DATA_BITWIDTH'b0000000100001001,
                    `W_DATA_BITWIDTH'b0000000100111100,
                    `W_DATA_BITWIDTH'b0000000101100110,
                    `W_DATA_BITWIDTH'b0000000101100101,
                    `W_DATA_BITWIDTH'b1111111000010001,
                    `W_DATA_BITWIDTH'b0000000110110101,
                    `W_DATA_BITWIDTH'b0000001000001111,
                    `W_DATA_BITWIDTH'b0000000111011010,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b1111111100001000,
                    `W_DATA_BITWIDTH'b0000000010001110,
                    `W_DATA_BITWIDTH'b1111111011101111,
                    `W_DATA_BITWIDTH'b1111111011001101,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b0000000101010000,
                    `W_DATA_BITWIDTH'b0000000101010000
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
                '{
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111111100100001,
                    `W_DATA_BITWIDTH'b1111111011010011,
                    `W_DATA_BITWIDTH'b1111111010000100,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b1111111011111100,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111111001011101,
                    `W_DATA_BITWIDTH'b1111111100010101,
                    `W_DATA_BITWIDTH'b1111111101010011,
                    `W_DATA_BITWIDTH'b1111111100000110,
                    `W_DATA_BITWIDTH'b1111111001111001,
                    `W_DATA_BITWIDTH'b1111111101100110,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b1111111010000001,
                    `W_DATA_BITWIDTH'b0000000011111001,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b1111111100100010,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b0000000010110010,
                    `W_DATA_BITWIDTH'b1111111101100101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b0000000100100110,
                    `W_DATA_BITWIDTH'b0000000010111100,
                    `W_DATA_BITWIDTH'b1111111101100101,
                    `W_DATA_BITWIDTH'b1111111010111001,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b1111111100001100,
                    `W_DATA_BITWIDTH'b1111111010011111,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b0000000011001011,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b0000000011010100,
                    `W_DATA_BITWIDTH'b0000000010000101,
                    `W_DATA_BITWIDTH'b0000000011111010,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b0000000010010001,
                    `W_DATA_BITWIDTH'b0000000011010010,
                    `W_DATA_BITWIDTH'b0000000010010100,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b0000000011111010,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b0000000100111100,
                    `W_DATA_BITWIDTH'b1111111101010101,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111101000111,
                    `W_DATA_BITWIDTH'b0000000011111010,
                    `W_DATA_BITWIDTH'b0000000011000001,
                    `W_DATA_BITWIDTH'b0000000101000101,
                    `W_DATA_BITWIDTH'b1111111011010000,
                    `W_DATA_BITWIDTH'b1111111001101011,
                    `W_DATA_BITWIDTH'b1111111010100111,
                    `W_DATA_BITWIDTH'b1111111011010001,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000110101011,
                    `W_DATA_BITWIDTH'b0000000011011010,
                    `W_DATA_BITWIDTH'b0000000100010010,
                    `W_DATA_BITWIDTH'b0000000101000000,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000100111011,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b1111111010100001,
                    `W_DATA_BITWIDTH'b0000000101000010,
                    `W_DATA_BITWIDTH'b1111111011101001,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111111010110110,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b1111111010010010,
                    `W_DATA_BITWIDTH'b0000000011111001,
                    `W_DATA_BITWIDTH'b0000000011111001,
                    `W_DATA_BITWIDTH'b1111111001111101,
                    `W_DATA_BITWIDTH'b0000000011101000,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000101011110,
                    `W_DATA_BITWIDTH'b1111110111101100,
                    `W_DATA_BITWIDTH'b0000000110101001,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000100110111,
                    `W_DATA_BITWIDTH'b1111110100110000,
                    `W_DATA_BITWIDTH'b0000000110000111,
                    `W_DATA_BITWIDTH'b1111111011100010,
                    `W_DATA_BITWIDTH'b1111111010000110,
                    `W_DATA_BITWIDTH'b1111111001000001,
                    `W_DATA_BITWIDTH'b1111110100100101,
                    `W_DATA_BITWIDTH'b1111111100101100,
                    `W_DATA_BITWIDTH'b1111111001000111,
                    `W_DATA_BITWIDTH'b0000000011010110,
                    `W_DATA_BITWIDTH'b0000000110101010,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111100000111,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b1111111000001100,
                    `W_DATA_BITWIDTH'b0000000101100111,
                    `W_DATA_BITWIDTH'b0000000111111010,
                    `W_DATA_BITWIDTH'b0000000111010110,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b0000000101001011,
                    `W_DATA_BITWIDTH'b0000000111111000,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b0000000101001000,
                    `W_DATA_BITWIDTH'b1111110100110011,
                    `W_DATA_BITWIDTH'b0000000110100100,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111111011001001,
                    `W_DATA_BITWIDTH'b0000001001110111,
                    `W_DATA_BITWIDTH'b0000001001011010,
                    `W_DATA_BITWIDTH'b0000000011001001,
                    `W_DATA_BITWIDTH'b1111111011101100,
                    `W_DATA_BITWIDTH'b1111111001110110,
                    `W_DATA_BITWIDTH'b0000000010000101,
                    `W_DATA_BITWIDTH'b1111111000101001,
                    `W_DATA_BITWIDTH'b1111111001100101,
                    `W_DATA_BITWIDTH'b0000000101101010,
                    `W_DATA_BITWIDTH'b1111111100111010,
                    `W_DATA_BITWIDTH'b1111111001001101,
                    `W_DATA_BITWIDTH'b1111111101011101,
                    `W_DATA_BITWIDTH'b0000000011010111,
                    `W_DATA_BITWIDTH'b1111110111000101,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111101111111,
                    `W_DATA_BITWIDTH'b1111111100111001,
                    `W_DATA_BITWIDTH'b1111111011100011,
                    `W_DATA_BITWIDTH'b1111111101001001,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011010010,
                    `W_DATA_BITWIDTH'b1111111100100100,
                    `W_DATA_BITWIDTH'b1111111011110000,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b0000000011110010,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111000110011,
                    `W_DATA_BITWIDTH'b0000000101110101,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b0000000010101001,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b1111111100110111,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b0000000100100110,
                    `W_DATA_BITWIDTH'b1111111000010011,
                    `W_DATA_BITWIDTH'b1111111100001001,
                    `W_DATA_BITWIDTH'b1111111101000001,
                    `W_DATA_BITWIDTH'b1111111100011111,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b1111111101101101,
                    `W_DATA_BITWIDTH'b1111111100011010,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000100110011,
                    `W_DATA_BITWIDTH'b0000000100010110,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b1111111100110101,
                    `W_DATA_BITWIDTH'b0000000010101001,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111011000010,
                    `W_DATA_BITWIDTH'b0000000010010101,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b0000000010001000,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b0000000011001010,
                    `W_DATA_BITWIDTH'b1111111101001001,
                    `W_DATA_BITWIDTH'b0000000011010011,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111111100001000,
                    `W_DATA_BITWIDTH'b1111111011010111,
                    `W_DATA_BITWIDTH'b0000000011100001,
                    `W_DATA_BITWIDTH'b0000000101110111,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b1111111011010101,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b0000000010000101,
                    `W_DATA_BITWIDTH'b0000000101110001,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000100001110,
                    `W_DATA_BITWIDTH'b1111111011000010,
                    `W_DATA_BITWIDTH'b1111111011100100,
                    `W_DATA_BITWIDTH'b1111111101110100,
                    `W_DATA_BITWIDTH'b1111111101101110,
                    `W_DATA_BITWIDTH'b1111111101001000,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111101010010,
                    `W_DATA_BITWIDTH'b1111111001110010,
                    `W_DATA_BITWIDTH'b0000000010100000,
                    `W_DATA_BITWIDTH'b1111111100011100,
                    `W_DATA_BITWIDTH'b0000000011110110,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b0000000010101001,
                    `W_DATA_BITWIDTH'b1111111100010110,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b1111111001010000,
                    `W_DATA_BITWIDTH'b1111111011111111,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b1111111011100011,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b1111111100110100,
                    `W_DATA_BITWIDTH'b1111111010110010,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111111100010111,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000011010010,
                    `W_DATA_BITWIDTH'b0000000110010010,
                    `W_DATA_BITWIDTH'b0000000011110101,
                    `W_DATA_BITWIDTH'b1111111101010110,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b0000000100000100,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b0000000111101000,
                    `W_DATA_BITWIDTH'b0000001000111011,
                    `W_DATA_BITWIDTH'b0000000111010000,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b1111111101100000,
                    `W_DATA_BITWIDTH'b0000000101100011,
                    `W_DATA_BITWIDTH'b1111110110110001,
                    `W_DATA_BITWIDTH'b0000001000011111,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b1111111000011100,
                    `W_DATA_BITWIDTH'b0000000111110101,
                    `W_DATA_BITWIDTH'b1111111100110000,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b1111110110101110,
                    `W_DATA_BITWIDTH'b0000000101000001,
                    `W_DATA_BITWIDTH'b0000000110100011,
                    `W_DATA_BITWIDTH'b0000000100111011,
                    `W_DATA_BITWIDTH'b0000000100001000,
                    `W_DATA_BITWIDTH'b1111110101001010,
                    `W_DATA_BITWIDTH'b1111111000101010,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111100110000,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111110111010001,
                    `W_DATA_BITWIDTH'b1111111101000111,
                    `W_DATA_BITWIDTH'b0000000011110100,
                    `W_DATA_BITWIDTH'b0000000110101110,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000100100111,
                    `W_DATA_BITWIDTH'b1111110111010011,
                    `W_DATA_BITWIDTH'b0000000110101101,
                    `W_DATA_BITWIDTH'b0000000011010110,
                    `W_DATA_BITWIDTH'b0000000101110110,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b0000000011100000,
                    `W_DATA_BITWIDTH'b1111111100111110,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b1111111101101111,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b0000000011011101,
                    `W_DATA_BITWIDTH'b1111111100000011,
                    `W_DATA_BITWIDTH'b1111111011101111,
                    `W_DATA_BITWIDTH'b0000000011011101,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111101010010,
                    `W_DATA_BITWIDTH'b1111111010010101,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b0000000010101111,
                    `W_DATA_BITWIDTH'b0000000110111111,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b1111111101100000,
                    `W_DATA_BITWIDTH'b1111111100011101,
                    `W_DATA_BITWIDTH'b0000001000011001,
                    `W_DATA_BITWIDTH'b1111111010001010,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b1111111100101100,
                    `W_DATA_BITWIDTH'b1111111001110110,
                    `W_DATA_BITWIDTH'b0000000011111101,
                    `W_DATA_BITWIDTH'b0000000100110101,
                    `W_DATA_BITWIDTH'b1111111000111011,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000011010110,
                    `W_DATA_BITWIDTH'b1111111011101111,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111010010011,
                    `W_DATA_BITWIDTH'b1111111100111010,
                    `W_DATA_BITWIDTH'b1111111011111110,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b1111111100001001,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b0000000010011010,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b1111111001110100,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b0000000100110101,
                    `W_DATA_BITWIDTH'b1111111011010100,
                    `W_DATA_BITWIDTH'b0000001000110110,
                    `W_DATA_BITWIDTH'b0000000101100111,
                    `W_DATA_BITWIDTH'b0000000101010011,
                    `W_DATA_BITWIDTH'b1111111001110111,
                    `W_DATA_BITWIDTH'b1111111101000001,
                    `W_DATA_BITWIDTH'b0000000101111101,
                    `W_DATA_BITWIDTH'b1111111010000100,
                    `W_DATA_BITWIDTH'b0000000110011110,
                    `W_DATA_BITWIDTH'b0000000101010101,
                    `W_DATA_BITWIDTH'b0000000100100000,
                    `W_DATA_BITWIDTH'b1111111010100000,
                    `W_DATA_BITWIDTH'b1111110110011101,
                    `W_DATA_BITWIDTH'b1111111101000001,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b1111111100000101,
                    `W_DATA_BITWIDTH'b1111110010111001,
                    `W_DATA_BITWIDTH'b0000001000011100,
                    `W_DATA_BITWIDTH'b0000000010110110,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b1111110010011011,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111110101111011,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b0000000111010110,
                    `W_DATA_BITWIDTH'b1111111100100001,
                    `W_DATA_BITWIDTH'b1111111000100001,
                    `W_DATA_BITWIDTH'b1111111001011001,
                    `W_DATA_BITWIDTH'b1111111010111100,
                    `W_DATA_BITWIDTH'b1111111000101001,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111001000101,
                    `W_DATA_BITWIDTH'b0000000010010010,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111101001000,
                    `W_DATA_BITWIDTH'b1111111101101010,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b1111111011000001,
                    `W_DATA_BITWIDTH'b1111111010110011,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b0000000100011011,
                    `W_DATA_BITWIDTH'b1111111000110110,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111111000010011,
                    `W_DATA_BITWIDTH'b1111111100100101,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b0000000110010110,
                    `W_DATA_BITWIDTH'b0000000010110101,
                    `W_DATA_BITWIDTH'b1111111101001011,
                    `W_DATA_BITWIDTH'b1111111101010100,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b1111111101100100,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111111100101110,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111111001100011,
                    `W_DATA_BITWIDTH'b0000000110011110,
                    `W_DATA_BITWIDTH'b0000000101110111,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b1111111101101111,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000100101111,
                    `W_DATA_BITWIDTH'b1111111101100001,
                    `W_DATA_BITWIDTH'b0000000101110000,
                    `W_DATA_BITWIDTH'b0000000101010010,
                    `W_DATA_BITWIDTH'b0000000110000111,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000100111110,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b1111111010110101,
                    `W_DATA_BITWIDTH'b1111111101111011,
                    `W_DATA_BITWIDTH'b0000000100010101,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b0000000100001011,
                    `W_DATA_BITWIDTH'b0000000010001001,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000100000001,
                    `W_DATA_BITWIDTH'b0000000100111111,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b0000000010110001,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111110110110000,
                    `W_DATA_BITWIDTH'b1111111101000011,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b0000000010101010,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b0000000011001101,
                    `W_DATA_BITWIDTH'b0000000100100110,
                    `W_DATA_BITWIDTH'b1111111101110000,
                    `W_DATA_BITWIDTH'b1111111100110010,
                    `W_DATA_BITWIDTH'b0000000010010101,
                    `W_DATA_BITWIDTH'b0000000101010110,
                    `W_DATA_BITWIDTH'b0000000011011000,
                    `W_DATA_BITWIDTH'b0000000010111101,
                    `W_DATA_BITWIDTH'b0000000010110100,
                    `W_DATA_BITWIDTH'b0000000011100010,
                    `W_DATA_BITWIDTH'b1111111101110100,
                    `W_DATA_BITWIDTH'b0000000010101101,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b0000000100100010,
                    `W_DATA_BITWIDTH'b0000000011010111,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111100000101,
                    `W_DATA_BITWIDTH'b1111110110010000,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b1111111011111011,
                    `W_DATA_BITWIDTH'b1111111011100001,
                    `W_DATA_BITWIDTH'b0000000101011000,
                    `W_DATA_BITWIDTH'b0000000010000001,
                    `W_DATA_BITWIDTH'b0000000011011000,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b1111110110101100,
                    `W_DATA_BITWIDTH'b1111111100010110,
                    `W_DATA_BITWIDTH'b1111111100001100,
                    `W_DATA_BITWIDTH'b1111111100100101,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b0000000010111010,
                    `W_DATA_BITWIDTH'b1111111010001110,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b1111111000010010,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b1111111010001110,
                    `W_DATA_BITWIDTH'b1111111010110101,
                    `W_DATA_BITWIDTH'b0000000010111111,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111100000101,
                    `W_DATA_BITWIDTH'b1111111000000110,
                    `W_DATA_BITWIDTH'b1111111101100010,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b0000000100100010,
                    `W_DATA_BITWIDTH'b0000000110000001,
                    `W_DATA_BITWIDTH'b0000000100000000,
                    `W_DATA_BITWIDTH'b0000001001000010,
                    `W_DATA_BITWIDTH'b0000001001000010
                };
                localparam logic signed [`W_DATA_BITWIDTH-1:0] w_data_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
                '{
                    `W_DATA_BITWIDTH'b0000000010100010,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b1111111011000000,
                    `W_DATA_BITWIDTH'b1111111101100100,
                    `W_DATA_BITWIDTH'b0000000011010001,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b0000000011010100,
                    `W_DATA_BITWIDTH'b1111111011110100,
                    `W_DATA_BITWIDTH'b1111111010010100,
                    `W_DATA_BITWIDTH'b0000000010010010,
                    `W_DATA_BITWIDTH'b1111111001110100,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b0000000011000111,
                    `W_DATA_BITWIDTH'b1111111100111010,
                    `W_DATA_BITWIDTH'b1111111101110111,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b1111111100011011,
                    `W_DATA_BITWIDTH'b0000000100110101,
                    `W_DATA_BITWIDTH'b1111111011111001,
                    `W_DATA_BITWIDTH'b1111111100000010,
                    `W_DATA_BITWIDTH'b0000000101001111,
                    `W_DATA_BITWIDTH'b1111111101011000,
                    `W_DATA_BITWIDTH'b0000000100000010,
                    `W_DATA_BITWIDTH'b1111111100101010,
                    `W_DATA_BITWIDTH'b1111111011001011,
                    `W_DATA_BITWIDTH'b1111111100100110,
                    `W_DATA_BITWIDTH'b0000000010010000,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b1111111011111100,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b1111111101110101,
                    `W_DATA_BITWIDTH'b0000000100101100,
                    `W_DATA_BITWIDTH'b0000000010101010,
                    `W_DATA_BITWIDTH'b0000000100101011,
                    `W_DATA_BITWIDTH'b1111111101010011,
                    `W_DATA_BITWIDTH'b1111111101100011,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b1111111010110010,
                    `W_DATA_BITWIDTH'b1111111010000100,
                    `W_DATA_BITWIDTH'b1111111101000110,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b0000000101000111,
                    `W_DATA_BITWIDTH'b0000001000110101,
                    `W_DATA_BITWIDTH'b1111111010010101,
                    `W_DATA_BITWIDTH'b0000000010010110,
                    `W_DATA_BITWIDTH'b0000000011111111,
                    `W_DATA_BITWIDTH'b0000000011100110,
                    `W_DATA_BITWIDTH'b1111111010000101,
                    `W_DATA_BITWIDTH'b0000000010101100,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111101110001,
                    `W_DATA_BITWIDTH'b0000000011100111,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b0000000011011010,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b0000000100010000,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b0000000011111100,
                    `W_DATA_BITWIDTH'b0000000011101100,
                    `W_DATA_BITWIDTH'b0000000100011001,
                    `W_DATA_BITWIDTH'b1111111000101110,
                    `W_DATA_BITWIDTH'b0000000111111110,
                    `W_DATA_BITWIDTH'b1111111001111000,
                    `W_DATA_BITWIDTH'b1111111100110011,
                    `W_DATA_BITWIDTH'b1111111000101101,
                    `W_DATA_BITWIDTH'b0000000011000011,
                    `W_DATA_BITWIDTH'b1111110111100011,
                    `W_DATA_BITWIDTH'b1111111011001111,
                    `W_DATA_BITWIDTH'b0000001011111010,
                    `W_DATA_BITWIDTH'b0000000100011000,
                    `W_DATA_BITWIDTH'b0000000110000001,
                    `W_DATA_BITWIDTH'b1111111011100101,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b1111110111100100,
                    `W_DATA_BITWIDTH'b1111111101111010,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b0000000101101110,
                    `W_DATA_BITWIDTH'b0000000011111110,
                    `W_DATA_BITWIDTH'b0000001000101110,
                    `W_DATA_BITWIDTH'b1111111000011001,
                    `W_DATA_BITWIDTH'b0000000100000001,
                    `W_DATA_BITWIDTH'b0000000101010111,
                    `W_DATA_BITWIDTH'b1111111001001100,
                    `W_DATA_BITWIDTH'b1111111011111101,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000110101010,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b1111111001011101,
                    `W_DATA_BITWIDTH'b1111111100001100,
                    `W_DATA_BITWIDTH'b0000000010101010,
                    `W_DATA_BITWIDTH'b1111110110110001,
                    `W_DATA_BITWIDTH'b1111111101101101,
                    `W_DATA_BITWIDTH'b1111110110111000,
                    `W_DATA_BITWIDTH'b0000001010000111,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b0000000100100111,
                    `W_DATA_BITWIDTH'b0000000100000001,
                    `W_DATA_BITWIDTH'b1111110110111110,
                    `W_DATA_BITWIDTH'b0000000110101001,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b1111110100100011,
                    `W_DATA_BITWIDTH'b0000000011101100,
                    `W_DATA_BITWIDTH'b1111111000000111,
                    `W_DATA_BITWIDTH'b1111111100001011,
                    `W_DATA_BITWIDTH'b1111111011010000,
                    `W_DATA_BITWIDTH'b1111111001000101,
                    `W_DATA_BITWIDTH'b1111111101011111,
                    `W_DATA_BITWIDTH'b1111110110100000,
                    `W_DATA_BITWIDTH'b1111111001111111,
                    `W_DATA_BITWIDTH'b0000000101101110,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b1111111001111010,
                    `W_DATA_BITWIDTH'b0000000010100111,
                    `W_DATA_BITWIDTH'b0000000100010011,
                    `W_DATA_BITWIDTH'b1111111011010001,
                    `W_DATA_BITWIDTH'b0000000101010111,
                    `W_DATA_BITWIDTH'b1111111010111000,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b1111111100010111,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b0000000010011011,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b1111111100111101,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b0000000011111111,
                    `W_DATA_BITWIDTH'b0000000101011001,
                    `W_DATA_BITWIDTH'b0000000011010100,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b1111111101011001,
                    `W_DATA_BITWIDTH'b0000000010011000,
                    `W_DATA_BITWIDTH'b1111111010001001,
                    `W_DATA_BITWIDTH'b0000000100000111,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b0000000010011001,
                    `W_DATA_BITWIDTH'b1111111100010011,
                    `W_DATA_BITWIDTH'b1111111001111111,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111011100000,
                    `W_DATA_BITWIDTH'b0000000101111010,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111001111010,
                    `W_DATA_BITWIDTH'b0000000011101100,
                    `W_DATA_BITWIDTH'b1111111011001000,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000011000101,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000011001000,
                    `W_DATA_BITWIDTH'b1111111001100100,
                    `W_DATA_BITWIDTH'b0000000100100000,
                    `W_DATA_BITWIDTH'b1111111101010000,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b1111111011110010,
                    `W_DATA_BITWIDTH'b1111110111010100,
                    `W_DATA_BITWIDTH'b1111111011101101,
                    `W_DATA_BITWIDTH'b1111111011001010,
                    `W_DATA_BITWIDTH'b1111111001101101,
                    `W_DATA_BITWIDTH'b1111111101110010,
                    `W_DATA_BITWIDTH'b1111111100010000,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000010011101,
                    `W_DATA_BITWIDTH'b0000000100000101,
                    `W_DATA_BITWIDTH'b1111111100001110,
                    `W_DATA_BITWIDTH'b0000000100111000,
                    `W_DATA_BITWIDTH'b1111111001111100,
                    `W_DATA_BITWIDTH'b1111111101010011,
                    `W_DATA_BITWIDTH'b1111111100101000,
                    `W_DATA_BITWIDTH'b1111111100010001,
                    `W_DATA_BITWIDTH'b0000000011011111,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111101011010,
                    `W_DATA_BITWIDTH'b1111110111101111,
                    `W_DATA_BITWIDTH'b1111111100111111,
                    `W_DATA_BITWIDTH'b1111111100111101,
                    `W_DATA_BITWIDTH'b0000000010100001,
                    `W_DATA_BITWIDTH'b0000000100100011,
                    `W_DATA_BITWIDTH'b0000000010010011,
                    `W_DATA_BITWIDTH'b1111110110101010,
                    `W_DATA_BITWIDTH'b1111111010011000,
                    `W_DATA_BITWIDTH'b0000000010000100,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b1111111100100111,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111001111101,
                    `W_DATA_BITWIDTH'b1111111011011101,
                    `W_DATA_BITWIDTH'b1111111010101100,
                    `W_DATA_BITWIDTH'b0000000010001000,
                    `W_DATA_BITWIDTH'b1111111000110010,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b1111111011110101,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000100111010,
                    `W_DATA_BITWIDTH'b1111111011001001,
                    `W_DATA_BITWIDTH'b0000000011111000,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b1111111011011011,
                    `W_DATA_BITWIDTH'b1111111011000010,
                    `W_DATA_BITWIDTH'b1111111010111111,
                    `W_DATA_BITWIDTH'b1111111011101100,
                    `W_DATA_BITWIDTH'b0000000010001111,
                    `W_DATA_BITWIDTH'b1111111010011101,
                    `W_DATA_BITWIDTH'b1111111101111101,
                    `W_DATA_BITWIDTH'b0000000011101110,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b0000000011000001,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b1111111101001110,
                    `W_DATA_BITWIDTH'b1111111010110011,
                    `W_DATA_BITWIDTH'b0000000101001100,
                    `W_DATA_BITWIDTH'b1111111010101000,
                    `W_DATA_BITWIDTH'b1111111011110011,
                    `W_DATA_BITWIDTH'b1111111000011101,
                    `W_DATA_BITWIDTH'b0000000010001101,
                    `W_DATA_BITWIDTH'b1111111010100100,
                    `W_DATA_BITWIDTH'b0000000010000010,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b1111111100111000,
                    `W_DATA_BITWIDTH'b0000000101100101,
                    `W_DATA_BITWIDTH'b0000000101000110,
                    `W_DATA_BITWIDTH'b1111111011011100,
                    `W_DATA_BITWIDTH'b0000000010011111,
                    `W_DATA_BITWIDTH'b1111111000110101,
                    `W_DATA_BITWIDTH'b0000000100100111,
                    `W_DATA_BITWIDTH'b1111110010101100,
                    `W_DATA_BITWIDTH'b1111110101111001,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b1111111010010111,
                    `W_DATA_BITWIDTH'b1111111001100101,
                    `W_DATA_BITWIDTH'b0000000101010110,
                    `W_DATA_BITWIDTH'b0000000010011001,
                    `W_DATA_BITWIDTH'b0000001010001010,
                    `W_DATA_BITWIDTH'b1111111000111101,
                    `W_DATA_BITWIDTH'b0000000011110011,
                    `W_DATA_BITWIDTH'b1111111001000111,
                    `W_DATA_BITWIDTH'b1111111010100111,
                    `W_DATA_BITWIDTH'b1111111000110000,
                    `W_DATA_BITWIDTH'b1111111000101011,
                    `W_DATA_BITWIDTH'b0000000100100000,
                    `W_DATA_BITWIDTH'b0000000011011011,
                    `W_DATA_BITWIDTH'b1111111100111011,
                    `W_DATA_BITWIDTH'b0000000010001011,
                    `W_DATA_BITWIDTH'b0000000111001010,
                    `W_DATA_BITWIDTH'b0000000101001000,
                    `W_DATA_BITWIDTH'b1111111001011001,
                    `W_DATA_BITWIDTH'b0000000101011010,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111111101111110,
                    `W_DATA_BITWIDTH'b1111111010101010,
                    `W_DATA_BITWIDTH'b0000000011110000,
                    `W_DATA_BITWIDTH'b1111111100101011,
                    `W_DATA_BITWIDTH'b0000000010100110,
                    `W_DATA_BITWIDTH'b1111111100111101,
                    `W_DATA_BITWIDTH'b0000000100001100,
                    `W_DATA_BITWIDTH'b0000000101000100,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b0000000011001010,
                    `W_DATA_BITWIDTH'b1111111011110010,
                    `W_DATA_BITWIDTH'b1111111011101011,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000100001011,
                    `W_DATA_BITWIDTH'b0000000011110000,
                    `W_DATA_BITWIDTH'b1111111011000011,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b0000000100011101,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111111101111000,
                    `W_DATA_BITWIDTH'b0000000101010111,
                    `W_DATA_BITWIDTH'b0000000010010001,
                    `W_DATA_BITWIDTH'b1111111101011110,
                    `W_DATA_BITWIDTH'b0000000110110001,
                    `W_DATA_BITWIDTH'b0000000100011111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b0000001000001001,
                    `W_DATA_BITWIDTH'b0000000010011010,
                    `W_DATA_BITWIDTH'b0000000100011010,
                    `W_DATA_BITWIDTH'b0000000110010110,
                    `W_DATA_BITWIDTH'b0000000010011110,
                    `W_DATA_BITWIDTH'b0000000110111000,
                    `W_DATA_BITWIDTH'b0000000011111101,
                    `W_DATA_BITWIDTH'b1111111001011110,
                    `W_DATA_BITWIDTH'b0000000011111011,
                    `W_DATA_BITWIDTH'b1111111100010100,
                    `W_DATA_BITWIDTH'b0000000011101101,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b0000000011010101,
                    `W_DATA_BITWIDTH'b1111111100111001,
                    `W_DATA_BITWIDTH'b0000000010100000,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b1111110111110110,
                    `W_DATA_BITWIDTH'b0000000101110100,
                    `W_DATA_BITWIDTH'b0000000110001101,
                    `W_DATA_BITWIDTH'b1111111001110000,
                    `W_DATA_BITWIDTH'b1111111100101111,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b0000000010001110,
                    `W_DATA_BITWIDTH'b0000000101110011,
                    `W_DATA_BITWIDTH'b1111111101100111,
                    `W_DATA_BITWIDTH'b1111110101111011,
                    `W_DATA_BITWIDTH'b0000001001101010,
                    `W_DATA_BITWIDTH'b0000000100110000,
                    `W_DATA_BITWIDTH'b1111110001100010,
                    `W_DATA_BITWIDTH'b0000001001110100,
                    `W_DATA_BITWIDTH'b0000000111000100,
                    `W_DATA_BITWIDTH'b1111111011110111,
                    `W_DATA_BITWIDTH'b1111110110100111,
                    `W_DATA_BITWIDTH'b0000000011101011,
                    `W_DATA_BITWIDTH'b1111111000001000,
                    `W_DATA_BITWIDTH'b1111111101001000,
                    `W_DATA_BITWIDTH'b0000000110011101,
                    `W_DATA_BITWIDTH'b1111111010011010,
                    `W_DATA_BITWIDTH'b1111110100100100,
                    `W_DATA_BITWIDTH'b0000000101000100,
                    `W_DATA_BITWIDTH'b0000000110101011,
                    `W_DATA_BITWIDTH'b1111111010111010,
                    `W_DATA_BITWIDTH'b1111111101101000,
                    `W_DATA_BITWIDTH'b1111111101011100,
                    `W_DATA_BITWIDTH'b0000000100010111,
                    `W_DATA_BITWIDTH'b0000000101100010,
                    `W_DATA_BITWIDTH'b1111111000011100,
                    `W_DATA_BITWIDTH'b0000000011001011,
                    `W_DATA_BITWIDTH'b1111111100000011,
                    `W_DATA_BITWIDTH'b1111111011010111,
                    `W_DATA_BITWIDTH'b0000000101111110,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b1111110011111000,
                    `W_DATA_BITWIDTH'b1111111001001011,
                    `W_DATA_BITWIDTH'b0000000010100101,
                    `W_DATA_BITWIDTH'b1111111011100011,
                    `W_DATA_BITWIDTH'b1111111001001100,
                    `W_DATA_BITWIDTH'b1111111100011000,
                    `W_DATA_BITWIDTH'b1111111001110010,
                    `W_DATA_BITWIDTH'b1111111101110100,
                    `W_DATA_BITWIDTH'b0000000101101000,
                    `W_DATA_BITWIDTH'b1111111001101100,
                    `W_DATA_BITWIDTH'b1111111010110000,
                    `W_DATA_BITWIDTH'b1111111101111001,
                    `W_DATA_BITWIDTH'b0000000011111011,
                    `W_DATA_BITWIDTH'b1111111010010100,
                    `W_DATA_BITWIDTH'b0000000101010000,
                    `W_DATA_BITWIDTH'b1111111100001010,
                    `W_DATA_BITWIDTH'b1111111011110001,
                    `W_DATA_BITWIDTH'b0000000011101010,
                    `W_DATA_BITWIDTH'b1111111101011011,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b1111111000101000,
                    `W_DATA_BITWIDTH'b1111111100111100,
                    `W_DATA_BITWIDTH'b0000000101001000,
                    `W_DATA_BITWIDTH'b0000000110000010,
                    `W_DATA_BITWIDTH'b1111111010110001,
                    `W_DATA_BITWIDTH'b0000000010110101,
                    `W_DATA_BITWIDTH'b1111111001011100,
                    `W_DATA_BITWIDTH'b0000000011001110,
                    `W_DATA_BITWIDTH'b1111111100010101,
                    `W_DATA_BITWIDTH'b1111111101001101,
                    `W_DATA_BITWIDTH'b1111111011011111,
                    `W_DATA_BITWIDTH'b0000000011110111,
                    `W_DATA_BITWIDTH'b1111111010101110,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b1111111100100010,
                    `W_DATA_BITWIDTH'b0000000011100100,
                    `W_DATA_BITWIDTH'b0000000100001000,
                    `W_DATA_BITWIDTH'b1111111100100000,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000101000101,
                    `W_DATA_BITWIDTH'b0000000011000001,
                    `W_DATA_BITWIDTH'b0000000010101110,
                    `W_DATA_BITWIDTH'b1111111100101101,
                    `W_DATA_BITWIDTH'b1111111011111111,
                    `W_DATA_BITWIDTH'b0000000011101001,
                    `W_DATA_BITWIDTH'b0000000010111100,
                    `W_DATA_BITWIDTH'b0000000010101011,
                    `W_DATA_BITWIDTH'b0000000011011100,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b0000000010010111,
                    `W_DATA_BITWIDTH'b0000000100101011,
                    `W_DATA_BITWIDTH'b0000000101101101,
                    `W_DATA_BITWIDTH'b1111111101110110,
                    `W_DATA_BITWIDTH'b1111110101001100,
                    `W_DATA_BITWIDTH'b1111111100100011,
                    `W_DATA_BITWIDTH'b1111111101000101,
                    `W_DATA_BITWIDTH'b0000000010100011,
                    `W_DATA_BITWIDTH'b1111111101010111,
                    `W_DATA_BITWIDTH'b1111111011111101,
                    `W_DATA_BITWIDTH'b1111111011111010,
                    `W_DATA_BITWIDTH'b0000000100101111,
                    `W_DATA_BITWIDTH'b0000000010000011,
                    `W_DATA_BITWIDTH'b0000000011101111,
                    `W_DATA_BITWIDTH'b0000000010001100,
                    `W_DATA_BITWIDTH'b0000000010001110,
                    `W_DATA_BITWIDTH'b1111111101100001,
                    `W_DATA_BITWIDTH'b0000000010000110,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b0000000010111011,
                    `W_DATA_BITWIDTH'b0000000010110000,
                    `W_DATA_BITWIDTH'b0000000100000111,
                    `W_DATA_BITWIDTH'b0000000100001111,
                    `W_DATA_BITWIDTH'b1111111011000001,
                    `W_DATA_BITWIDTH'b1111111001100000,
                    `W_DATA_BITWIDTH'b1111111100110110,
                    `W_DATA_BITWIDTH'b1111110110000111,
                    `W_DATA_BITWIDTH'b1111111100101001,
                    `W_DATA_BITWIDTH'b1111111010011101,
                    `W_DATA_BITWIDTH'b0000000101000110,
                    `W_DATA_BITWIDTH'b0000000101100011,
                    `W_DATA_BITWIDTH'b0000000010100101,
                    `W_DATA_BITWIDTH'b0000000101011011,
                    `W_DATA_BITWIDTH'b1111111100011111,
                    `W_DATA_BITWIDTH'b1111111001100010,
                    `W_DATA_BITWIDTH'b0000000100011000,
                    `W_DATA_BITWIDTH'b0000000100010011,
                    `W_DATA_BITWIDTH'b1111111101110011,
                    `W_DATA_BITWIDTH'b0000000011001100,
                    `W_DATA_BITWIDTH'b0000000100111011,
                    `W_DATA_BITWIDTH'b1111111010001011,
                    `W_DATA_BITWIDTH'b1111111100000111,
                    `W_DATA_BITWIDTH'b0000001001000101,
                    `W_DATA_BITWIDTH'b1111111101001111,
                    `W_DATA_BITWIDTH'b1111111010010110,
                    `W_DATA_BITWIDTH'b0000001000111001,
                    `W_DATA_BITWIDTH'b0000000111110000,
                    `W_DATA_BITWIDTH'b1111111101101001,
                    `W_DATA_BITWIDTH'b1111111001101010,
                    `W_DATA_BITWIDTH'b1111111011001000,
                    `W_DATA_BITWIDTH'b0000000011011011,
                    `W_DATA_BITWIDTH'b1111110110110101,
                    `W_DATA_BITWIDTH'b1111111100000000,
                    `W_DATA_BITWIDTH'b0000000010101000,
                    `W_DATA_BITWIDTH'b0000000100000110,
                    `W_DATA_BITWIDTH'b0000001000000111,
                    `W_DATA_BITWIDTH'b0000000100111100,
                    `W_DATA_BITWIDTH'b0000000100111100
                };

            // w_c_idx
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s0 [0:`W_C_LENGTH_L1_S0-1] =
                '{
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s1 [0:`W_C_LENGTH_L1_S1-1] =
                '{
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l1_s2 [0:`W_C_LENGTH_L1_S2-1] =
                '{
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00001
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s0 [0:`W_C_LENGTH_L2_S0-1] =
                '{
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01110
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s1 [0:`W_C_LENGTH_L2_S1-1] =
                '{
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01110
                };
                localparam logic [`W_C_BITWIDTH-1:0] w_c_idx_l2_s2 [0:`W_C_LENGTH_L2_S2-1] =
                '{
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01001,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01100,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00001,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00110,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01111,
                    `W_C_BITWIDTH'b00000,
                    `W_C_BITWIDTH'b00010,
                    `W_C_BITWIDTH'b00011,
                    `W_C_BITWIDTH'b00100,
                    `W_C_BITWIDTH'b00101,
                    `W_C_BITWIDTH'b00111,
                    `W_C_BITWIDTH'b01000,
                    `W_C_BITWIDTH'b01010,
                    `W_C_BITWIDTH'b01011,
                    `W_C_BITWIDTH'b01101,
                    `W_C_BITWIDTH'b01110,
                    `W_C_BITWIDTH'b01110
                };

            // w_r_idx
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };
                localparam logic [`W_R_BITWIDTH-1:0] w_r_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
                '{
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b10,
                    `W_R_BITWIDTH'b00,
                    `W_R_BITWIDTH'b01,
                    `W_R_BITWIDTH'b01
                };

            // w_k_idx
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };
                localparam logic [`W_K_BITWIDTH-1:0] w_k_idx_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
                '{
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00000,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00001,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00010,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00011,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00100,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00101,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00110,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b00111,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01000,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01001,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01010,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01011,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01100,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01101,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01110,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111,
                    `W_K_BITWIDTH'b01111
                };

            // w_pos_ptr
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s0 [0:`W_R_LENGTH_L1_S0-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00000000000,
                    `W_POS_PTR_BITWIDTH'b00000000010,
                    `W_POS_PTR_BITWIDTH'b00000000100,
                    `W_POS_PTR_BITWIDTH'b00000000110,
                    `W_POS_PTR_BITWIDTH'b00000001000,
                    `W_POS_PTR_BITWIDTH'b00000001010,
                    `W_POS_PTR_BITWIDTH'b00000001101,
                    `W_POS_PTR_BITWIDTH'b00000010000,
                    `W_POS_PTR_BITWIDTH'b00000010011,
                    `W_POS_PTR_BITWIDTH'b00000010110,
                    `W_POS_PTR_BITWIDTH'b00000011001,
                    `W_POS_PTR_BITWIDTH'b00000011100,
                    `W_POS_PTR_BITWIDTH'b00000011110,
                    `W_POS_PTR_BITWIDTH'b00000100000,
                    `W_POS_PTR_BITWIDTH'b00000100011,
                    `W_POS_PTR_BITWIDTH'b00000100110,
                    `W_POS_PTR_BITWIDTH'b00000101001,
                    `W_POS_PTR_BITWIDTH'b00000101100,
                    `W_POS_PTR_BITWIDTH'b00000101110,
                    `W_POS_PTR_BITWIDTH'b00000110000,
                    `W_POS_PTR_BITWIDTH'b00000110011,
                    `W_POS_PTR_BITWIDTH'b00000110101,
                    `W_POS_PTR_BITWIDTH'b00000111000,
                    `W_POS_PTR_BITWIDTH'b00000111010,
                    `W_POS_PTR_BITWIDTH'b00000111100,
                    `W_POS_PTR_BITWIDTH'b00000111111,
                    `W_POS_PTR_BITWIDTH'b00001000010,
                    `W_POS_PTR_BITWIDTH'b00001000100,
                    `W_POS_PTR_BITWIDTH'b00001000111,
                    `W_POS_PTR_BITWIDTH'b00001001010,
                    `W_POS_PTR_BITWIDTH'b00001001101,
                    `W_POS_PTR_BITWIDTH'b00001001110,
                    `W_POS_PTR_BITWIDTH'b00001010000,
                    `W_POS_PTR_BITWIDTH'b00001010010,
                    `W_POS_PTR_BITWIDTH'b00001010101,
                    `W_POS_PTR_BITWIDTH'b00001011000,
                    `W_POS_PTR_BITWIDTH'b00001011011,
                    `W_POS_PTR_BITWIDTH'b00001011110,
                    `W_POS_PTR_BITWIDTH'b00001100001,
                    `W_POS_PTR_BITWIDTH'b00001100100,
                    `W_POS_PTR_BITWIDTH'b00001100110,
                    `W_POS_PTR_BITWIDTH'b00001101000,
                    `W_POS_PTR_BITWIDTH'b00001101011,
                    `W_POS_PTR_BITWIDTH'b00001101101,
                    `W_POS_PTR_BITWIDTH'b00001110000,
                    `W_POS_PTR_BITWIDTH'b00001110010,
                    `W_POS_PTR_BITWIDTH'b00001110101,
                    `W_POS_PTR_BITWIDTH'b00001110101
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s1 [0:`W_R_LENGTH_L1_S1-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00001111011,
                    `W_POS_PTR_BITWIDTH'b00001111101,
                    `W_POS_PTR_BITWIDTH'b00001111111,
                    `W_POS_PTR_BITWIDTH'b00010000010,
                    `W_POS_PTR_BITWIDTH'b00010000101,
                    `W_POS_PTR_BITWIDTH'b00010001000,
                    `W_POS_PTR_BITWIDTH'b00010001011,
                    `W_POS_PTR_BITWIDTH'b00010001110,
                    `W_POS_PTR_BITWIDTH'b00010010001,
                    `W_POS_PTR_BITWIDTH'b00010010100,
                    `W_POS_PTR_BITWIDTH'b00010010111,
                    `W_POS_PTR_BITWIDTH'b00010011001,
                    `W_POS_PTR_BITWIDTH'b00010011100,
                    `W_POS_PTR_BITWIDTH'b00010011111,
                    `W_POS_PTR_BITWIDTH'b00010100010,
                    `W_POS_PTR_BITWIDTH'b00010100101,
                    `W_POS_PTR_BITWIDTH'b00010101000,
                    `W_POS_PTR_BITWIDTH'b00010101011,
                    `W_POS_PTR_BITWIDTH'b00010101110,
                    `W_POS_PTR_BITWIDTH'b00010110000,
                    `W_POS_PTR_BITWIDTH'b00010110010,
                    `W_POS_PTR_BITWIDTH'b00010110101,
                    `W_POS_PTR_BITWIDTH'b00010111000,
                    `W_POS_PTR_BITWIDTH'b00010111010,
                    `W_POS_PTR_BITWIDTH'b00010111101,
                    `W_POS_PTR_BITWIDTH'b00011000000,
                    `W_POS_PTR_BITWIDTH'b00011000011,
                    `W_POS_PTR_BITWIDTH'b00011000110,
                    `W_POS_PTR_BITWIDTH'b00011001001,
                    `W_POS_PTR_BITWIDTH'b00011001100,
                    `W_POS_PTR_BITWIDTH'b00011001110,
                    `W_POS_PTR_BITWIDTH'b00011010000,
                    `W_POS_PTR_BITWIDTH'b00011010010,
                    `W_POS_PTR_BITWIDTH'b00011010011,
                    `W_POS_PTR_BITWIDTH'b00011010110,
                    `W_POS_PTR_BITWIDTH'b00011011001,
                    `W_POS_PTR_BITWIDTH'b00011011100,
                    `W_POS_PTR_BITWIDTH'b00011011111,
                    `W_POS_PTR_BITWIDTH'b00011100010,
                    `W_POS_PTR_BITWIDTH'b00011100101,
                    `W_POS_PTR_BITWIDTH'b00011101000,
                    `W_POS_PTR_BITWIDTH'b00011101011,
                    `W_POS_PTR_BITWIDTH'b00011101110,
                    `W_POS_PTR_BITWIDTH'b00011110000,
                    `W_POS_PTR_BITWIDTH'b00011110010,
                    `W_POS_PTR_BITWIDTH'b00011110101,
                    `W_POS_PTR_BITWIDTH'b00011111000,
                    `W_POS_PTR_BITWIDTH'b00011111000
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l1_s2 [0:`W_R_LENGTH_L1_S2-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00011111101,
                    `W_POS_PTR_BITWIDTH'b00100000000,
                    `W_POS_PTR_BITWIDTH'b00100000010,
                    `W_POS_PTR_BITWIDTH'b00100000101,
                    `W_POS_PTR_BITWIDTH'b00100001000,
                    `W_POS_PTR_BITWIDTH'b00100001001,
                    `W_POS_PTR_BITWIDTH'b00100001100,
                    `W_POS_PTR_BITWIDTH'b00100001111,
                    `W_POS_PTR_BITWIDTH'b00100010010,
                    `W_POS_PTR_BITWIDTH'b00100010101,
                    `W_POS_PTR_BITWIDTH'b00100011000,
                    `W_POS_PTR_BITWIDTH'b00100011011,
                    `W_POS_PTR_BITWIDTH'b00100011110,
                    `W_POS_PTR_BITWIDTH'b00100100000,
                    `W_POS_PTR_BITWIDTH'b00100100011,
                    `W_POS_PTR_BITWIDTH'b00100100110,
                    `W_POS_PTR_BITWIDTH'b00100101000,
                    `W_POS_PTR_BITWIDTH'b00100101011,
                    `W_POS_PTR_BITWIDTH'b00100101110,
                    `W_POS_PTR_BITWIDTH'b00100110000,
                    `W_POS_PTR_BITWIDTH'b00100110011,
                    `W_POS_PTR_BITWIDTH'b00100110110,
                    `W_POS_PTR_BITWIDTH'b00100111000,
                    `W_POS_PTR_BITWIDTH'b00100111010,
                    `W_POS_PTR_BITWIDTH'b00100111101,
                    `W_POS_PTR_BITWIDTH'b00101000000,
                    `W_POS_PTR_BITWIDTH'b00101000011,
                    `W_POS_PTR_BITWIDTH'b00101000110,
                    `W_POS_PTR_BITWIDTH'b00101001001,
                    `W_POS_PTR_BITWIDTH'b00101001100,
                    `W_POS_PTR_BITWIDTH'b00101001111,
                    `W_POS_PTR_BITWIDTH'b00101010000,
                    `W_POS_PTR_BITWIDTH'b00101010001,
                    `W_POS_PTR_BITWIDTH'b00101010010,
                    `W_POS_PTR_BITWIDTH'b00101010100,
                    `W_POS_PTR_BITWIDTH'b00101010111,
                    `W_POS_PTR_BITWIDTH'b00101011010,
                    `W_POS_PTR_BITWIDTH'b00101011101,
                    `W_POS_PTR_BITWIDTH'b00101011111,
                    `W_POS_PTR_BITWIDTH'b00101100010,
                    `W_POS_PTR_BITWIDTH'b00101100100,
                    `W_POS_PTR_BITWIDTH'b00101100111,
                    `W_POS_PTR_BITWIDTH'b00101101010,
                    `W_POS_PTR_BITWIDTH'b00101101100,
                    `W_POS_PTR_BITWIDTH'b00101101110,
                    `W_POS_PTR_BITWIDTH'b00101110001,
                    `W_POS_PTR_BITWIDTH'b00101110100,
                    `W_POS_PTR_BITWIDTH'b00101110100
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s0 [0:`W_R_LENGTH_L2_S0-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00000000000,
                    `W_POS_PTR_BITWIDTH'b00000001010,
                    `W_POS_PTR_BITWIDTH'b00000010001,
                    `W_POS_PTR_BITWIDTH'b00000011001,
                    `W_POS_PTR_BITWIDTH'b00000011111,
                    `W_POS_PTR_BITWIDTH'b00000101001,
                    `W_POS_PTR_BITWIDTH'b00000110001,
                    `W_POS_PTR_BITWIDTH'b00000111001,
                    `W_POS_PTR_BITWIDTH'b00001000101,
                    `W_POS_PTR_BITWIDTH'b00001010001,
                    `W_POS_PTR_BITWIDTH'b00001011110,
                    `W_POS_PTR_BITWIDTH'b00001100110,
                    `W_POS_PTR_BITWIDTH'b00001110100,
                    `W_POS_PTR_BITWIDTH'b00001111111,
                    `W_POS_PTR_BITWIDTH'b00010001001,
                    `W_POS_PTR_BITWIDTH'b00010010100,
                    `W_POS_PTR_BITWIDTH'b00010011011,
                    `W_POS_PTR_BITWIDTH'b00010100101,
                    `W_POS_PTR_BITWIDTH'b00010101110,
                    `W_POS_PTR_BITWIDTH'b00010110101,
                    `W_POS_PTR_BITWIDTH'b00010111110,
                    `W_POS_PTR_BITWIDTH'b00011000100,
                    `W_POS_PTR_BITWIDTH'b00011001101,
                    `W_POS_PTR_BITWIDTH'b00011010110,
                    `W_POS_PTR_BITWIDTH'b00011100000,
                    `W_POS_PTR_BITWIDTH'b00011101011,
                    `W_POS_PTR_BITWIDTH'b00011111000,
                    `W_POS_PTR_BITWIDTH'b00100000110,
                    `W_POS_PTR_BITWIDTH'b00100010000,
                    `W_POS_PTR_BITWIDTH'b00100011001,
                    `W_POS_PTR_BITWIDTH'b00100011110,
                    `W_POS_PTR_BITWIDTH'b00100101001,
                    `W_POS_PTR_BITWIDTH'b00100110111,
                    `W_POS_PTR_BITWIDTH'b00101000000,
                    `W_POS_PTR_BITWIDTH'b00101001010,
                    `W_POS_PTR_BITWIDTH'b00101010100,
                    `W_POS_PTR_BITWIDTH'b00101100001,
                    `W_POS_PTR_BITWIDTH'b00101101101,
                    `W_POS_PTR_BITWIDTH'b00101110111,
                    `W_POS_PTR_BITWIDTH'b00110000011,
                    `W_POS_PTR_BITWIDTH'b00110001101,
                    `W_POS_PTR_BITWIDTH'b00110010110,
                    `W_POS_PTR_BITWIDTH'b00110011110,
                    `W_POS_PTR_BITWIDTH'b00110100101,
                    `W_POS_PTR_BITWIDTH'b00110101111,
                    `W_POS_PTR_BITWIDTH'b00110110110,
                    `W_POS_PTR_BITWIDTH'b00111000011,
                    `W_POS_PTR_BITWIDTH'b00111000011
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s1 [0:`W_R_LENGTH_L2_S1-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b00111011010,
                    `W_POS_PTR_BITWIDTH'b00111100100,
                    `W_POS_PTR_BITWIDTH'b00111101110,
                    `W_POS_PTR_BITWIDTH'b00111110111,
                    `W_POS_PTR_BITWIDTH'b01000000000,
                    `W_POS_PTR_BITWIDTH'b01000001000,
                    `W_POS_PTR_BITWIDTH'b01000001110,
                    `W_POS_PTR_BITWIDTH'b01000011000,
                    `W_POS_PTR_BITWIDTH'b01000011110,
                    `W_POS_PTR_BITWIDTH'b01000101010,
                    `W_POS_PTR_BITWIDTH'b01000110101,
                    `W_POS_PTR_BITWIDTH'b01001000010,
                    `W_POS_PTR_BITWIDTH'b01001001111,
                    `W_POS_PTR_BITWIDTH'b01001011100,
                    `W_POS_PTR_BITWIDTH'b01001100001,
                    `W_POS_PTR_BITWIDTH'b01001101011,
                    `W_POS_PTR_BITWIDTH'b01001110100,
                    `W_POS_PTR_BITWIDTH'b01001111100,
                    `W_POS_PTR_BITWIDTH'b01010000100,
                    `W_POS_PTR_BITWIDTH'b01010001111,
                    `W_POS_PTR_BITWIDTH'b01010010111,
                    `W_POS_PTR_BITWIDTH'b01010011110,
                    `W_POS_PTR_BITWIDTH'b01010101010,
                    `W_POS_PTR_BITWIDTH'b01010110010,
                    `W_POS_PTR_BITWIDTH'b01010111110,
                    `W_POS_PTR_BITWIDTH'b01011001000,
                    `W_POS_PTR_BITWIDTH'b01011010101,
                    `W_POS_PTR_BITWIDTH'b01011100010,
                    `W_POS_PTR_BITWIDTH'b01011100111,
                    `W_POS_PTR_BITWIDTH'b01011101111,
                    `W_POS_PTR_BITWIDTH'b01011110100,
                    `W_POS_PTR_BITWIDTH'b01100000000,
                    `W_POS_PTR_BITWIDTH'b01100001000,
                    `W_POS_PTR_BITWIDTH'b01100010001,
                    `W_POS_PTR_BITWIDTH'b01100011011,
                    `W_POS_PTR_BITWIDTH'b01100100101,
                    `W_POS_PTR_BITWIDTH'b01100110100,
                    `W_POS_PTR_BITWIDTH'b01100111111,
                    `W_POS_PTR_BITWIDTH'b01101001000,
                    `W_POS_PTR_BITWIDTH'b01101010011,
                    `W_POS_PTR_BITWIDTH'b01101011111,
                    `W_POS_PTR_BITWIDTH'b01101100111,
                    `W_POS_PTR_BITWIDTH'b01101101101,
                    `W_POS_PTR_BITWIDTH'b01101110111,
                    `W_POS_PTR_BITWIDTH'b01101111110,
                    `W_POS_PTR_BITWIDTH'b01110000101,
                    `W_POS_PTR_BITWIDTH'b01110010001,
                    `W_POS_PTR_BITWIDTH'b01110010001
                };
                localparam logic [`W_POS_PTR_BITWIDTH-1:0] w_pos_ptr_l2_s2 [0:`W_R_LENGTH_L2_S2-1] =
                '{
                    `W_POS_PTR_BITWIDTH'b01110100110,
                    `W_POS_PTR_BITWIDTH'b01110101100,
                    `W_POS_PTR_BITWIDTH'b01110110011,
                    `W_POS_PTR_BITWIDTH'b01110111011,
                    `W_POS_PTR_BITWIDTH'b01111000011,
                    `W_POS_PTR_BITWIDTH'b01111001011,
                    `W_POS_PTR_BITWIDTH'b01111010010,
                    `W_POS_PTR_BITWIDTH'b01111011110,
                    `W_POS_PTR_BITWIDTH'b01111100111,
                    `W_POS_PTR_BITWIDTH'b01111110001,
                    `W_POS_PTR_BITWIDTH'b01111111101,
                    `W_POS_PTR_BITWIDTH'b10000001001,
                    `W_POS_PTR_BITWIDTH'b10000010101,
                    `W_POS_PTR_BITWIDTH'b10000011111,
                    `W_POS_PTR_BITWIDTH'b10000100111,
                    `W_POS_PTR_BITWIDTH'b10000110100,
                    `W_POS_PTR_BITWIDTH'b10000111100,
                    `W_POS_PTR_BITWIDTH'b10001000110,
                    `W_POS_PTR_BITWIDTH'b10001001110,
                    `W_POS_PTR_BITWIDTH'b10001010100,
                    `W_POS_PTR_BITWIDTH'b10001100001,
                    `W_POS_PTR_BITWIDTH'b10001101100,
                    `W_POS_PTR_BITWIDTH'b10001110111,
                    `W_POS_PTR_BITWIDTH'b10010000000,
                    `W_POS_PTR_BITWIDTH'b10010000110,
                    `W_POS_PTR_BITWIDTH'b10010010001,
                    `W_POS_PTR_BITWIDTH'b10010011011,
                    `W_POS_PTR_BITWIDTH'b10010101001,
                    `W_POS_PTR_BITWIDTH'b10010110010,
                    `W_POS_PTR_BITWIDTH'b10010111000,
                    `W_POS_PTR_BITWIDTH'b10011000000,
                    `W_POS_PTR_BITWIDTH'b10011001011,
                    `W_POS_PTR_BITWIDTH'b10011010100,
                    `W_POS_PTR_BITWIDTH'b10011011100,
                    `W_POS_PTR_BITWIDTH'b10011101100,
                    `W_POS_PTR_BITWIDTH'b10011110111,
                    `W_POS_PTR_BITWIDTH'b10100000011,
                    `W_POS_PTR_BITWIDTH'b10100001100,
                    `W_POS_PTR_BITWIDTH'b10100010101,
                    `W_POS_PTR_BITWIDTH'b10100011110,
                    `W_POS_PTR_BITWIDTH'b10100100011,
                    `W_POS_PTR_BITWIDTH'b10100101100,
                    `W_POS_PTR_BITWIDTH'b10100110100,
                    `W_POS_PTR_BITWIDTH'b10100111011,
                    `W_POS_PTR_BITWIDTH'b10100111111,
                    `W_POS_PTR_BITWIDTH'b10101000001,
                    `W_POS_PTR_BITWIDTH'b10101001101,
                    `W_POS_PTR_BITWIDTH'b10101001101
                };



    // ========================== Logic (Wire) =============================================
        // ----------------------- For PE ------- unfinished------------------------
            logic                                  i_start_PEs;
            // IA bundle
            logic        [$clog2(`IA_ROW)-1:0]     i_ia_h;
            logic        [$clog2(`IA_COL)-1:0]     i_ia_w;
            logic signed [`IA_DATA_BITWIDTH-1:0]   i_ia_data   [0:`IA_CHANNEL-1];
            logic        [`IA_C_BITWIDTH-1:0]      i_ia_c_idx  [0:`IA_CHANNEL-1];
            logic        [$clog2(`IA_CHANNEL)-1:0] i_ia_iters; // ---------------------- need discussion -> 0
            logic        [$clog2(`IA_CHANNEL)-1:0] i_ia_len;
            // W bundle
            logic        [1:0]                     i_w_s;
            logic signed [`W_DATA_BITWIDTH-1:0]    i_w_data    [0:`W_C_LENGTH-1]; 
            logic        [`W_C_BITWIDTH-1:0]       i_w_c_idx   [0:`W_C_LENGTH-1];
            logic        [`W_POS_PTR_BITWIDTH-1:0] i_pos_ptr   [0:`W_R_LENGTH-1];
            logic        [`W_R_BITWIDTH-1:0]       i_r_idx     [0:`W_R_LENGTH-1];
            logic        [`W_K_BITWIDTH-1:0]       i_k_idx     [0:`W_R_LENGTH-1];
            logic        [$clog2(`W_C_LENGTH)-1:0] i_w_iters;  // ---------------------- need discussion -> ceil(w_len/32)
            logic        [$clog2(`W_C_LENGTH)-1:0] i_w_len;
            // Output
            logic                                  o_finish_PE;
            logic signed [`IA_DATA_BITWIDTH-1:0]   o_OA        [0:`IA_ROW-1][0:`IA_CHANNEL-1];

	PE_TEMP pe_temp0(
        .i_rst_n        (rst),
		.i_clk          (clk),
        .i_start        (i_start_PEs),
        // IA bundle
        .i_ia_h         (i_ia_h),
        .i_ia_w         (i_ia_w),
        .i_ia_data      (i_ia_data),
        .i_ia_c_idx     (i_ia_c_idx ),
        .i_ia_iters     (i_ia_iters),
        .i_ia_len       (i_ia_len),
        // W bundle
        .i_w_s          (i_w_s),
        .i_w_data       (i_w_data),
        .i_w_c_idx      (i_w_c_idx),
        .i_pos_ptr      (i_pos_ptr),
        .i_r_idx        (i_r_idx),
        .i_k_idx        (i_k_idx),
        .i_w_iters      (i_w_iters),
        .i_w_len        (i_w_len),
        // Output
        .o_finish       (o_finish),
        .o_OA           (o_OA)
	);

	initial begin
		$fsdbDumpfile("pe_temp.fsdb");
		$fsdbDumpvars;
		$fsdbDumpMDA();
        // reset 
		rst = 1'b0;
		#(2*CLK)
		rst = 1'b1;

        for (int i = 0; i < 10; i++) @(posedge clk);




        for (int i = 0; i < 5000; i++) begin
            @(posedge clk);
            //-----------------------
                i_start_PEs = 1;
                // IA bundle
                i_ia_h      = 0;
                i_ia_w      = 0;
                for (int k=0; k < `IA_CHANNEL; k++) begin 
                    i_ia_data[k]  = (k<3) ? (2*k+1) : -2;
                    i_ia_c_idx[k] = (k<3) ? (k*k)  : 0;
                end
                i_ia_iters  = 0; // fixed
                i_ia_len    = 3;

                // W bundle
                i_w_s       = 0;
                for (int k=0; k < `W_C_LENGTH; k++) i_w_data[k]    = (k<`W_C_LENGTH_L1_S0) ? w_data_l1_s0[k]    : -1;
                for (int k=0; k < `W_C_LENGTH; k++) i_w_c_idx[k]   = (k<`W_C_LENGTH_L1_S0) ? w_c_idx_l1_s0[k]   : 0; 
                for (int k=0; k < `W_R_LENGTH; k++) i_pos_ptr[k]   = (k<`W_R_LENGTH_L1_S0) ? w_pos_ptr_l1_s0[k] : 0; 
                for (int k=0; k < `W_R_LENGTH; k++) i_r_idx[k]     = (k<`W_R_LENGTH_L1_S0) ? w_r_idx_l1_s0[k]   : 0; 
                for (int k=0; k < `W_R_LENGTH; k++) i_k_idx[k]     = (k<`W_R_LENGTH_L1_S0) ? w_k_idx_l1_s0[k]   : 0; 
                i_w_iters   = (`W_C_LENGTH_L1_S0 >> 5);
                i_w_len     = `W_C_LENGTH_L1_S0;

        end




        $finish;
    end
	initial begin
		#(50000*CLK)
		$display(".A.B.O.R.T.");
		$finish;
	end

endmodule
